* SPICE3 file created from gf180mcu_voidwalkers_sc_sdffrnq_4_flattened.ext - technology: gf180mcuD

.option scale=5n

.subckt gf180mcu_voidwalkers_sc_sdffrnq_4_flattened_pex VDD VSS A B S CLK RN Q
X0 a_n870_270# RN.t0 VDD.t4 VDD.t3 pfet_03v3 ad=51n pd=0.98m as=37.4n ps=0.9m w=340 l=60
X1 a_2090_270# S.t0 A.t1 VDD.t25 pfet_03v3 ad=22.1n pd=0.47m as=41.14n ps=0.922m w=340 l=60
X2 a_n1490_270# a_n1300_270# VSS.t29 VSS.t28 nfet_03v3 ad=21.93n pd=0.598m as=11.05n ps=0.3m w=170 l=60
X3 a_n1300_270# a_n870_270# VSS.t17 VSS.t16 nfet_03v3 ad=11.05n pd=0.3m as=18.7n ps=0.56m w=170 l=60
X4 a_120_270# a_n870_270# VSS.t15 VSS.t14 nfet_03v3 ad=11.05n pd=0.3m as=18.7n ps=0.56m w=170 l=60
X5 a_1370_270# CLK.t0 a_1620_320# VSS.t21 nfet_03v3 ad=11.05n pd=0.3m as=7.65n ps=0.26m w=170 l=60
X6 a_n730_520# CLK.t1 a_n430_810# VDD.t18 pfet_03v3 ad=22.1n pd=0.47m as=15.3n ps=0.43m w=340 l=60
X7 a_n340_270# CLK.t2 VSS.t20 VSS.t19 nfet_03v3 ad=30.6n pd=0.7m as=11.05n ps=0.3m w=170 l=60
X8 VDD.t1 a_n730_520# a_n780_810# VDD.t0 pfet_03v3 ad=30.6n pd=0.52m as=8.5n ps=0.39m w=340 l=60
X9 a_1620_810# a_120_270# VDD.t11 VDD.t10 pfet_03v3 ad=15.3n pd=0.43m as=22.1n ps=0.47m w=340 l=60
X10 a_2910_160# S.t1 VDD.t6 VDD.t5 pfet_03v3 ad=37.4n pd=0.9m as=44.2n ps=0.94m w=340 l=60
X11 a_2090_270# a_2910_160# A.t0 VSS.t2 nfet_03v3 ad=11.05n pd=0.3m as=20.57n ps=0.582m w=170 l=60
X12 VDD.t9 a_120_270# a_n90_810# VDD.t8 pfet_03v3 ad=22.1n pd=0.47m as=35.7n ps=0.55m w=340 l=60
X13 a_1710_650# CLK.t3 VDD.t20 VDD.t19 pfet_03v3 ad=61.2n pd=1.04m as=22.1n ps=0.47m w=340 l=60
X14 a_1270_810# a_n870_270# a_120_270# VDD.t16 pfet_03v3 ad=17n pd=0.44m as=37.4n ps=0.9m w=340 l=60
X15 a_n730_520# a_n340_270# a_n430_320# VSS.t5 nfet_03v3 ad=24.65n pd=0.46m as=7.65n ps=0.26m w=170 l=60
X16 a_1620_320# a_120_270# VSS.t9 VSS.t8 nfet_03v3 ad=7.65n pd=0.26m as=11.05n ps=0.3m w=170 l=60
X17 a_2910_160# S.t2 VSS.t24 VSS.t23 nfet_03v3 ad=18.7n pd=0.56m as=22.1n ps=0.6m w=170 l=60
X18 VSS.t1 a_n730_520# a_n1300_270# VSS.t0 nfet_03v3 ad=11.05n pd=0.3m as=11.05n ps=0.3m w=170 l=60
X19 B.t0 a_2910_160# a_2090_270# VDD.t2 pfet_03v3 ad=44.2n pd=0.94m as=22.1n ps=0.47m w=340 l=60
X20 a_70_320# CLK.t4 a_n730_520# VSS.t25 nfet_03v3 ad=4.25n pd=0.22m as=24.65n ps=0.46m w=170 l=60
X21 VDD.t29 a_n1490_270# Q.t0 VDD.t28 pfet_03v3 ad=22.1n pd=0.47m as=37.4n ps=0.9m w=340 l=60
X22 a_n90_810# a_n340_270# a_n730_520# VDD.t7 pfet_03v3 ad=35.7n pd=0.55m as=22.1n ps=0.47m w=340 l=60
X23 VSS.t7 a_120_270# a_70_320# VSS.t6 nfet_03v3 ad=11.05n pd=0.3m as=4.25n ps=0.22m w=170 l=60
X24 a_n430_810# a_n1300_270# VDD.t24 VDD.t23 pfet_03v3 ad=15.3n pd=0.43m as=30.6n ps=0.52m w=340 l=60
X25 VDD.t31 a_1370_270# a_1270_810# VDD.t30 pfet_03v3 ad=22.1n pd=0.47m as=17n ps=0.44m w=340 l=60
X26 a_1960_810# CLK.t5 a_1370_270# VDD.t14 pfet_03v3 ad=22.1n pd=0.47m as=22.1n ps=0.47m w=340 l=60
X27 a_1710_650# CLK.t6 VSS.t13 VSS.t12 nfet_03v3 ad=30.6n pd=0.7m as=11.05n ps=0.3m w=170 l=60
X28 a_n780_810# a_n870_270# a_n1300_270# VDD.t15 pfet_03v3 ad=8.5n pd=0.39m as=37.4n ps=0.9m w=340 l=60
X29 B.t1 S.t3 a_2090_270# VSS.t22 nfet_03v3 ad=22.1n pd=0.6m as=11.05n ps=0.3m w=170 l=60
X30 VDD.t13 a_2090_270# a_1960_810# VDD.t12 pfet_03v3 ad=22.1n pd=0.47m as=22.1n ps=0.47m w=340 l=60
X31 VSS.t31 a_n1490_270# Q.t1 VSS.t30 nfet_03v3 ad=11.05n pd=0.3m as=18.7n ps=0.56m w=170 l=60
X32 VSS.t33 a_1370_270# a_120_270# VSS.t32 nfet_03v3 ad=11.05n pd=0.3m as=11.05n ps=0.3m w=170 l=60
X33 a_1960_320# a_1710_650# a_1370_270# VSS.t18 nfet_03v3 ad=11.05n pd=0.3m as=11.05n ps=0.3m w=170 l=60
X34 a_n430_320# a_n1300_270# VSS.t27 VSS.t26 nfet_03v3 ad=7.65n pd=0.26m as=11.05n ps=0.3m w=170 l=60
X35 a_n1490_270# a_n1300_270# VDD.t22 VDD.t21 pfet_03v3 ad=43.86n pd=0.938m as=22.1n ps=0.47m w=340 l=60
X36 a_1370_270# a_1710_650# a_1620_810# VDD.t17 pfet_03v3 ad=22.1n pd=0.47m as=15.3n ps=0.43m w=340 l=60
X37 VSS.t11 a_2090_270# a_1960_320# VSS.t10 nfet_03v3 ad=11.05n pd=0.3m as=11.05n ps=0.3m w=170 l=60
X38 a_n870_270# RN.t1 VSS.t4 VSS.t3 nfet_03v3 ad=25.5n pd=0.64m as=18.7n ps=0.56m w=170 l=60
X39 a_n340_270# CLK.t7 VDD.t27 VDD.t26 pfet_03v3 ad=61.2n pd=1.04m as=22.1n ps=0.47m w=340 l=60
C0 a_120_270# a_n870_270# 0.74762f
C1 VDD a_n730_520# 0.67699f
C2 VDD a_1270_810# 0.00447f
C3 Q a_n1300_270# 0.00445f
C4 a_n340_270# RN 0.04143f
C5 B VDD 0.07746f
C6 a_120_270# a_1620_810# 0
C7 a_1960_810# a_1370_270# 0.01518f
C8 VDD a_1370_270# 0.87978f
C9 a_n430_810# a_n730_520# 0.0266f
C10 S A 0.01847f
C11 CLK RN 0.03174f
C12 VDD a_n780_810# 0.0075f
C13 RN a_n870_270# 0.10161f
C14 S a_2090_270# 0.07571f
C15 RN a_120_270# 0.07609f
C16 VDD a_1710_650# 0.24742f
C17 a_1960_810# a_1710_650# 0.00909f
C18 a_1620_320# a_120_270# 0.00243f
C19 VDD a_2910_160# 1.24042f
C20 VDD a_n340_270# 0.19764f
C21 B a_2090_270# 0.34499f
C22 a_2090_270# a_1370_270# 0.02911f
C23 CLK VDD 1.09472f
C24 a_n1300_270# a_n730_520# 0.63309f
C25 a_n90_810# a_n730_520# 0.012f
C26 a_n1490_270# a_n870_270# 0.00218f
C27 A a_1710_650# 0.07531f
C28 VDD a_n870_270# 1.65825f
C29 CLK a_n430_810# 0.00481f
C30 B S 0.05446f
C31 A a_2910_160# 0.01056f
C32 a_n780_810# a_n1300_270# 0.00967f
C33 VDD a_120_270# 1.61783f
C34 CLK A 0.03677f
C35 a_2090_270# a_1710_650# 0.63962f
C36 a_2090_270# a_2910_160# 0.0342f
C37 a_n430_810# a_120_270# 0
C38 a_n780_810# a_n730_520# 0.00338f
C39 S a_1710_650# 0
C40 CLK a_2090_270# 0.16066f
C41 S a_2910_160# 0.4729f
C42 VDD RN 0.19951f
C43 a_n340_270# a_n1300_270# 0.0224f
C44 a_n340_270# a_n90_810# 0.00286f
C45 CLK a_n1300_270# 0.03156f
C46 CLK a_n90_810# 0.03152f
C47 CLK S 0.00834f
C48 a_70_320# a_n730_520# 0.00163f
C49 a_n340_270# a_n730_520# 0.0914f
C50 a_n1300_270# a_n870_270# 0.10345f
C51 a_1710_650# a_1370_270# 0.188f
C52 B a_2910_160# 0.45603f
C53 a_2910_160# a_1370_270# 0
C54 a_1960_320# a_1370_270# 0.00759f
C55 CLK a_n730_520# 0.34176f
C56 a_n1300_270# a_120_270# 0
C57 a_n90_810# a_120_270# 0.00506f
C58 a_n730_520# a_n870_270# 0.11752f
C59 CLK a_1370_270# 0.05158f
C60 VDD a_n1490_270# 0.40639f
C61 a_1960_810# VDD 0.02719f
C62 RN a_2090_270# 0
C63 a_n870_270# a_1370_270# 0.04501f
C64 a_120_270# a_n730_520# 0.00704f
C65 a_120_270# a_1270_810# 0.02752f
C66 a_2910_160# a_1710_650# 0
C67 a_1960_320# a_1710_650# 0.0079f
C68 a_1620_810# a_1370_270# 0.02857f
C69 a_n430_320# a_n730_520# 0.01223f
C70 a_120_270# a_1370_270# 0.55679f
C71 Q a_n1490_270# 0.17056f
C72 Q VDD 0.23146f
C73 a_70_320# a_n340_270# 0.00429f
C74 CLK a_1710_650# 0.25807f
C75 VDD A 0.03946f
C76 CLK a_2910_160# 0.00499f
C77 RN a_n730_520# 0
C78 CLK a_n340_270# 0.55128f
C79 a_n340_270# a_n870_270# 0.03884f
C80 RN a_1370_270# 0
C81 VDD a_2090_270# 1.16453f
C82 a_120_270# a_1710_650# 0.03483f
C83 a_1620_320# a_1370_270# 0.00628f
C84 CLK a_n870_270# 0.06033f
C85 a_n340_270# a_120_270# 0.42613f
C86 a_n1300_270# a_n1490_270# 0.6795f
C87 VDD a_n1300_270# 0.67224f
C88 VDD a_n90_810# 0.0258f
C89 S VDD 0.4527f
C90 CLK a_120_270# 0.48194f
C91 a_n430_320# a_n340_270# 0
C92 A a_2090_270# 0.34378f
R0 RN.n0 RN.t0 32.8505
R1 RN.n0 RN.t1 24.9422
R2 RN RN.n0 8.0455
R3 VDD.t2 VDD.t5 666.668
R4 VDD.t21 VDD.t15 638.889
R5 VDD.n11 VDD.t25 625
R6 VDD.t3 VDD.t16 583.333
R7 VDD.t26 VDD.n12 458.334
R8 VDD.t7 VDD.t8 375
R9 VDD.t0 VDD.t23 333.334
R10 VDD.t25 VDD.t2 263.889
R11 VDD.t12 VDD.t19 263.889
R12 VDD.t14 VDD.t12 263.889
R13 VDD.t17 VDD.t14 263.889
R14 VDD.t30 VDD.t10 263.889
R15 VDD.t8 VDD.t26 263.889
R16 VDD.t18 VDD.t7 263.889
R17 VDD.t28 VDD.t21 263.889
R18 VDD.t19 VDD.n11 250
R19 VDD.t16 VDD.t30 222.222
R20 VDD.t10 VDD.t17 208.333
R21 VDD.n12 VDD.t3 208.333
R22 VDD.t23 VDD.t18 208.333
R23 VDD.t15 VDD.t0 152.779
R24 VDD.n13 VDD.t28 95.9338
R25 VDD.n12 VDD.n0 12.6005
R26 VDD.n6 VDD.t4 11.1026
R27 VDD.n11 VDD.n10 6.3005
R28 VDD.n15 VDD.n2 5.40621
R29 VDD.n16 VDD.n1 5.40621
R30 VDD.n10 VDD.t6 4.86098
R31 VDD.n8 VDD.n5 2.86381
R32 VDD.n9 VDD.n4 2.86381
R33 VDD.n14 VDD.n3 2.85935
R34 VDD.n2 VDD.t24 1.95638
R35 VDD.n2 VDD.t1 1.7505
R36 VDD.n7 VDD 1.5755
R37 VDD.n5 VDD.t11 1.33874
R38 VDD.n5 VDD.t31 1.33874
R39 VDD.n4 VDD.t20 1.33874
R40 VDD.n4 VDD.t13 1.33874
R41 VDD.n3 VDD.t22 1.33874
R42 VDD.n3 VDD.t29 1.33874
R43 VDD.n1 VDD.t27 1.33874
R44 VDD.n1 VDD.t9 1.33874
R45 VDD VDD.n17 1.17981
R46 VDD.n16 VDD.n15 0.534071
R47 VDD.n15 VDD.n14 0.501929
R48 VDD.n8 VDD.n7 0.473
R49 VDD.n9 VDD.n8 0.463357
R50 VDD.n17 VDD.n16 0.222286
R51 VDD.n10 VDD.n9 0.177286
R52 VDD.n13 VDD 0.109786
R53 VDD.n14 VDD.n13 0.100143
R54 VDD.n17 VDD.n0 0.0418793
R55 VDD.n6 VDD.n0 0.0289483
R56 VDD.n7 VDD.n6 0.0186034
R57 S.n1 S.t0 57.1838
R58 S.n0 S.t1 41.3672
R59 S.n2 S.n1 31.7555
R60 S.n0 S.t2 16.4255
R61 S.n1 S.t3 16.4255
R62 S S.n2 8.0755
R63 S.n2 S.n0 3.2855
R64 A A.t0 8.85718
R65 A A.t1 6.96624
R66 VSS.t22 VSS.t23 2836.36
R67 VSS.t19 VSS.t3 2836.36
R68 VSS.n12 VSS.t2 2659.09
R69 VSS.t28 VSS.t16 2540.91
R70 VSS.t3 VSS.t14 2304.55
R71 VSS.t2 VSS.t22 1122.73
R72 VSS.t10 VSS.t12 1122.73
R73 VSS.t18 VSS.t10 1122.73
R74 VSS.t21 VSS.t18 1122.73
R75 VSS.t32 VSS.t8 1122.73
R76 VSS.t14 VSS.t32 1122.73
R77 VSS.t6 VSS.t19 1122.73
R78 VSS.n13 VSS.t25 1122.73
R79 VSS.t26 VSS.t0 1122.73
R80 VSS.t30 VSS.t28 1122.73
R81 VSS.t12 VSS.n12 1063.64
R82 VSS.n13 VSS.t5 945.456
R83 VSS.t8 VSS.t21 886.365
R84 VSS.t5 VSS.t26 886.365
R85 VSS.n19 VSS.t30 719.491
R86 VSS.t25 VSS.t6 650
R87 VSS.n18 VSS.t0 650
R88 VSS.t16 VSS.n18 472.728
R89 VSS.n11 VSS.t24 9.58039
R90 VSS.n8 VSS.t15 8.92147
R91 VSS.n7 VSS.t4 8.92147
R92 VSS.n16 VSS.t17 8.92147
R93 VSS.n10 VSS.n5 6.51264
R94 VSS.n9 VSS.n6 6.51264
R95 VSS.n1 VSS.n0 6.50965
R96 VSS.n15 VSS.n2 6.49979
R97 VSS.n4 VSS.n3 6.46764
R98 VSS.n12 VSS.n11 5.2005
R99 VSS.n14 VSS.n13 5.2005
R100 VSS.n18 VSS.n17 5.2005
R101 VSS.n5 VSS.t13 2.40932
R102 VSS.n5 VSS.t11 2.40932
R103 VSS.n6 VSS.t9 2.40932
R104 VSS.n6 VSS.t33 2.40932
R105 VSS.n3 VSS.t20 2.40932
R106 VSS.n3 VSS.t7 2.40932
R107 VSS.n2 VSS.t27 2.40932
R108 VSS.n2 VSS.t1 2.40932
R109 VSS.n0 VSS.t29 2.40932
R110 VSS.n0 VSS.t31 2.40932
R111 VSS.n10 VSS.n9 0.463357
R112 VSS.n7 VSS.n4 0.309071
R113 VSS.n16 VSS.n1 0.276929
R114 VSS.n15 VSS.n14 0.260857
R115 VSS.n14 VSS.n4 0.254429
R116 VSS.n8 VSS.n7 0.251214
R117 VSS.n9 VSS.n8 0.244786
R118 VSS.n11 VSS.n10 0.177286
R119 VSS.n19 VSS.n1 0.138714
R120 VSS.n17 VSS.n15 0.132286
R121 VSS.n17 VSS.n16 0.113
R122 VSS VSS.n19 0.0712143
R123 CLK.n1 CLK.n0 170.333
R124 CLK.t3 CLK.t5 111.933
R125 CLK.t6 CLK.n1 91.8588
R126 CLK.t4 CLK.t1 75.0038
R127 CLK.t2 CLK.t7 69.9588
R128 CLK.n0 CLK.t4 59.0088
R129 CLK CLK.n2 39.6788
R130 CLK.n2 CLK.t3 34.0672
R131 CLK.n2 CLK.t6 28.5922
R132 CLK.n1 CLK.t0 22.5088
R133 CLK.n0 CLK.t2 22.5088
R134 B B.t1 8.85718
R135 B B.t0 4.42383
R136 Q Q.t0 11.4292
R137 Q Q.t1 8.96004
C93 B VSS 0.06655f
C94 A VSS 0.10075f
C95 S VSS 0.74919f
C96 RN VSS 0.30296f
C97 Q VSS 0.29394f
C98 CLK VSS 2.74665f
C99 VDD VSS 12.7941f
C100 a_1960_320# VSS 0.01499f 
C101 a_1620_320# VSS 0.01063f 
C102 a_70_320# VSS 0.00445f
C103 a_1620_810# VSS 0 
C104 a_2910_160# VSS 1.39006f 
C105 a_2090_270# VSS 0.27786f 
C106 a_1710_650# VSS 0.5979f 
C107 a_1370_270# VSS 0.3449f
C108 a_120_270# VSS 0.76519f 
C109 a_n340_270# VSS 0.70374f 
C110 a_n730_520# VSS 0.5225f 
C111 a_n1300_270# VSS 0.91157f 
C112 a_n1490_270# VSS 0.59162f
C113 a_n870_270# VSS 1.1529f 
.ends

magic
tech gf180mcuD
magscale 1 10
timestamp 1756129822
<< nwell >>
rect -260 300 1510 1020
<< pwell >>
rect -260 -250 1510 300
<< nmos >>
rect -60 -30 0 140
rect 130 -30 190 140
rect 580 -30 640 140
rect 770 -30 830 140
rect 1250 -30 1310 140
<< pmos >>
rect -60 460 0 800
rect 130 460 190 800
rect 580 460 640 800
rect 770 460 830 800
rect 1250 460 1310 800
<< ndiff >>
rect -170 120 -60 140
rect -170 -10 -150 120
rect -100 -10 -60 120
rect -170 -30 -60 -10
rect 0 120 130 140
rect 0 -10 40 120
rect 90 -10 130 120
rect 0 -30 130 -10
rect 190 120 319 140
rect 190 -10 230 120
rect 280 -10 319 120
rect 190 -30 319 -10
rect 459 120 580 140
rect 459 -10 490 120
rect 540 -10 580 120
rect 459 -30 580 -10
rect 640 120 770 140
rect 640 -10 680 120
rect 730 -10 770 120
rect 640 -30 770 -10
rect 830 120 960 140
rect 830 -10 870 120
rect 920 -10 960 120
rect 1120 120 1250 140
rect 830 -30 960 -10
rect 1120 -10 1160 120
rect 1210 -10 1250 120
rect 1120 -30 1250 -10
rect 1310 120 1420 140
rect 1310 -10 1350 120
rect 1400 -10 1420 120
rect 1310 -30 1420 -10
<< pdiff >>
rect -170 780 -60 800
rect -170 660 -150 780
rect -100 660 -60 780
rect -170 460 -60 660
rect 0 780 130 800
rect 0 660 40 780
rect 90 660 130 780
rect 0 600 130 660
rect 0 480 40 600
rect 90 480 130 600
rect 0 460 130 480
rect 190 780 319 800
rect 190 660 230 780
rect 280 660 319 780
rect 190 600 319 660
rect 190 480 230 600
rect 280 480 319 600
rect 190 460 319 480
rect 459 600 580 800
rect 459 480 490 600
rect 540 480 580 600
rect 459 460 580 480
rect 640 780 770 800
rect 640 660 680 780
rect 730 660 770 780
rect 640 600 770 660
rect 640 480 680 600
rect 730 480 770 600
rect 640 460 770 480
rect 830 780 960 800
rect 830 660 870 780
rect 920 660 960 780
rect 1120 780 1250 800
rect 830 600 960 660
rect 830 480 870 600
rect 920 480 960 600
rect 830 460 960 480
rect 1120 660 1160 780
rect 1210 660 1250 780
rect 1120 600 1250 660
rect 1120 480 1160 600
rect 1210 480 1250 600
rect 1120 460 1250 480
rect 1310 780 1420 800
rect 1310 660 1350 780
rect 1400 660 1420 780
rect 1310 600 1420 660
rect 1310 480 1350 600
rect 1400 480 1420 600
rect 1310 460 1420 480
<< ndiffc >>
rect -150 -10 -100 120
rect 40 -10 90 120
rect 230 -10 280 120
rect 490 -10 540 120
rect 680 -10 730 120
rect 870 -10 920 120
rect 1160 -10 1210 120
rect 1350 -10 1400 120
<< pdiffc >>
rect -150 660 -100 780
rect 40 660 90 780
rect 40 480 90 600
rect 230 660 280 780
rect 230 480 280 600
rect 490 480 540 600
rect 680 660 730 780
rect 680 480 730 600
rect 870 660 920 780
rect 870 480 920 600
rect 1160 660 1210 780
rect 1160 480 1210 600
rect 1350 660 1400 780
rect 1350 480 1400 600
<< psubdiff >>
rect -220 -150 -80 -130
rect -220 -200 -200 -150
rect -100 -200 -80 -150
rect -220 -220 -80 -200
<< nsubdiff >>
rect -170 970 -70 990
rect -170 920 -150 970
rect -90 920 -70 970
rect -170 900 -70 920
<< psubdiffcont >>
rect -200 -200 -100 -150
<< nsubdiffcont >>
rect -150 920 -90 970
<< polysilicon >>
rect 770 850 1100 900
rect -60 800 0 850
rect 130 800 190 850
rect 580 800 640 850
rect 770 800 830 850
rect 1020 830 1100 850
rect 1020 719 1036 830
rect 1085 719 1100 830
rect 1250 800 1310 850
rect 1020 700 1100 719
rect -60 290 0 460
rect 130 410 190 460
rect 130 390 450 410
rect 130 330 340 390
rect 430 330 450 390
rect 130 310 450 330
rect 580 360 640 460
rect 770 410 830 460
rect -60 270 80 290
rect -60 210 -40 270
rect 60 210 80 270
rect -60 190 80 210
rect -60 140 0 190
rect 130 140 190 310
rect 580 300 830 360
rect 770 290 830 300
rect 1250 290 1310 460
rect 770 270 1310 290
rect 770 210 1180 270
rect 1290 210 1310 270
rect 770 190 1310 210
rect 580 140 640 190
rect 770 140 830 190
rect 1250 140 1310 190
rect 1020 50 1100 70
rect -60 -80 0 -30
rect 130 -80 190 -30
rect 580 -130 640 -30
rect 770 -80 830 -30
rect 1020 -61 1036 50
rect 1085 -61 1100 50
rect 1020 -130 1100 -61
rect 1250 -80 1310 -30
rect 580 -190 1100 -130
<< polycontact >>
rect 1036 719 1085 830
rect 340 330 430 390
rect -40 210 60 270
rect 1180 210 1290 270
rect 1036 -61 1085 50
<< metal1 >>
rect -260 970 1510 1020
rect -260 920 -150 970
rect -90 920 1510 970
rect -260 900 1510 920
rect -160 780 -90 800
rect -160 660 -150 780
rect -100 660 -90 780
rect -160 120 -90 660
rect 30 780 101 900
rect 1020 830 1100 850
rect 30 660 40 780
rect 90 660 101 780
rect 30 600 101 660
rect 30 480 40 600
rect 90 590 101 600
rect 220 780 290 800
rect 220 660 230 780
rect 280 660 290 780
rect 220 600 290 660
rect 90 480 100 590
rect 30 460 100 480
rect 220 480 230 600
rect 280 480 290 600
rect 220 290 290 480
rect 340 780 740 800
rect 340 670 680 780
rect 340 390 430 670
rect 670 660 680 670
rect 730 660 740 780
rect 340 310 430 330
rect 480 600 550 620
rect 480 480 490 600
rect 540 480 550 600
rect -40 270 290 290
rect 60 210 290 270
rect 480 260 550 480
rect -40 190 290 210
rect -160 -10 -150 120
rect -100 -10 -90 120
rect -160 -30 -90 -10
rect 30 120 101 144
rect 30 -10 40 120
rect 90 -10 101 120
rect 30 -130 101 -10
rect 220 120 290 190
rect 430 170 550 260
rect 220 -10 230 120
rect 280 -10 290 120
rect 220 -30 290 -10
rect 480 120 550 170
rect 480 -10 490 120
rect 540 -10 550 120
rect 480 -30 550 -10
rect 670 600 740 660
rect 670 480 680 600
rect 730 480 740 600
rect 670 120 740 480
rect 860 780 930 800
rect 860 660 870 780
rect 920 660 930 780
rect 860 600 930 660
rect 860 480 870 600
rect 920 480 930 600
rect 860 260 930 480
rect 810 170 930 260
rect 670 -10 680 120
rect 730 -10 740 120
rect 670 -30 740 -10
rect 860 120 930 170
rect 860 -10 870 120
rect 920 -10 930 120
rect 860 -30 930 -10
rect 1020 719 1036 830
rect 1085 719 1100 830
rect 1020 410 1100 719
rect 1150 780 1220 900
rect 1150 660 1160 780
rect 1210 660 1220 780
rect 1150 600 1220 660
rect 1150 480 1160 600
rect 1210 480 1220 600
rect 1150 460 1220 480
rect 1340 780 1450 800
rect 1340 660 1350 780
rect 1400 660 1450 780
rect 1340 600 1450 660
rect 1340 480 1350 600
rect 1400 480 1450 600
rect 1340 460 1450 480
rect 1390 410 1450 460
rect 1020 330 1450 410
rect 1020 50 1100 330
rect 1160 210 1180 270
rect 1290 210 1310 270
rect 1160 190 1310 210
rect 1390 140 1450 330
rect 1020 -61 1036 50
rect 1085 -61 1100 50
rect 1020 -80 1100 -61
rect 1150 120 1220 140
rect 1150 -10 1160 120
rect 1210 -10 1220 120
rect 1150 -130 1220 -10
rect 1340 120 1450 140
rect 1340 -10 1350 120
rect 1400 -10 1450 120
rect 1340 -30 1450 -10
rect -260 -150 1510 -130
rect -260 -200 -200 -150
rect -100 -200 1510 -150
rect -260 -250 1510 -200
<< labels >>
flabel metal1 s -160 200 -90 400 0 FreeSans 400 0 0 0 OUT
port 2 nsew
flabel metal1 s 1180 210 1290 270 0 FreeSans 400 0 0 0 SELECTOR
port 3 nsew
flabel metal1 s -260 900 1510 1020 0 FreeSans 400 0 0 0 VDD
port 6 nsew
flabel metal1 s -260 -250 1510 -130 0 FreeSans 400 0 0 0 VSS
port 8 nsew
flabel metal1 s 450 190 530 240 0 FreeSans 400 0 0 0 INPUT_2
port 9 nsew
flabel metal1 s 830 190 910 240 0 FreeSans 400 0 0 0 INPUT_1
port 10 nsew
<< end >>

  X �     �      (UNNAMED)  >A�7KƧ�9D�/��ZT �     �      pfet_03v3_6DGS6C        ,��΂������΂  R���  R���������΂����          ,���h�������h  R���  R����������h����          ,���N�������N  R����  R�����������N����          ,���4�������4  R����  R�����������4����          ,����������  R���  R��������������          ,��� �������   R���  R���������� ����          ,������������  R����  R����������������          ,������������  R���h  R���h������������          ,������������  R  N  R  N������������          ,  �����  �  R  4  R  4����  �����          ,  	~����  	~  R    R  ����  	~����          ,  d����  d  R     R   ����  d����          ,  J����  J  R  �  R  �����  J����          ,  0����  0  R  �  R  �����  0����          ,  !����  !  R  %�  R  %�����  !����          ,  &�����  &�  R  +�  R  +�����  &�����          ,  ,�����  ,�  R  1~  R  1~����  ,�����          ,���:�������:  .���f  .���f�������:����          ,��� �������   .���L  .���L������� ����          ,����������  .���2  .���2�����������          ,������������  .���  .���������������          ,������������  .����  .����������������          ,����������  .����  .���������������          ,����������  .����  .���������������          ,������������  .����  .����������������          ,���j�������j  .   �  .   ��������j����          ,  P����  P  .  |  .  |����  P����          ,  6����  6  .  b  .  b����  6����          ,  ����    .  H  .  H����  ����          ,  ����    .  .  .  .����  ����          ,  �����  �  .    .  ����  �����          ,  "�����  "�  .  #�  .  #�����  "�����          ,  (�����  (�  .  )�  .  )�����  (�����          ,  .�����  .�  .  /�  .  /�����  .�����      !    ,  ,  h  ,  D    D    h  ,  h      !    ,  �  h  �  D  �  D  �  h  �  h      !    ,    h    D  �  D  �  h    h      !    ,  	�  h  	�  D  
�  D  
�  h  	�  h      !    ,  �  h  �  D  �  D  �  h  �  h      !    ,  �  h  �  D  �  D  �  h  �  h      !    ,  �  h  �  D  �  D  �  h  �  h      !    ,  �  h  �  D  l  D  l  h  �  h      !    ,  �  h  �  D  �  D  �  h  �  h      !    ,  v  h  v  D  R  D  R  h  v  h      !    ,  �  h  �  D  �  D  �  h  �  h      !    ,  !\  h  !\  D  "8  D  "8  h  !\  h      !    ,  $�  h  $�  D  %l  D  %l  h  $�  h      !    ,  'B  h  'B  D  (  D  (  h  'B  h      !    ,  *v  h  *v  D  +R  D  +R  h  *v  h      !    ,  -(  h  -(  D  .  D  .  h  -(  h      !    ,  0\  h  0\  D  18  D  18  h  0\  h      !    ,  ,����  ,   n     n  ����  ,����      !    ,  �����  �   n  �   n  �����  �����      !    ,  ����     n  �   n  �����  ����      !    ,  	�����  	�   n  
�   n  
�����  	�����      !    ,  �����  �   n  �   n  �����  �����      !    ,  �����  �   n  �   n  �����  �����      !    ,  �����  �   n  �   n  �����  �����      !    ,  �����  �   n  l   n  l����  �����      !    ,  �����  �   n  �   n  �����  �����      !    ,  v����  v   n  R   n  R����  v����      !    ,  �����  �   n  �   n  �����  �����      !    ,  !\����  !\   n  "8   n  "8����  !\����      !    ,  $�����  $�   n  %l   n  %l����  $�����      !    ,  'B����  'B   n  (   n  (����  'B����      !    ,  *v����  *v   n  +R   n  +R����  *v����      !    ,  -(����  -(   n  .   n  .����  -(����      !    ,  0\����  0\   n  18   n  18����  0\����      !    ,  ,����  ,����  ����  ����  ,����      !    ,  �����  �����  �����  �����  �����      !    ,  ����  ����  �����  �����  ����      !    ,  	�����  	�����  
�����  
�����  	�����      !    ,  �����  �����  �����  �����  �����      !    ,  �����  �����  �����  �����  �����      !    ,  �����  �����  �����  �����  �����      !    ,  �����  �����  l����  l����  �����      !    ,  �����  �����  �����  �����  �����      !    ,  v����  v����  R����  R����  v����      !    ,  �����  �����  �����  �����  �����      !    ,  !\����  !\����  "8����  "8����  !\����      !    ,  $�����  $�����  %l����  %l����  $�����      !    ,  'B����  'B����  (����  (����  'B����      !    ,  *v����  *v����  +R����  +R����  *v����      !    ,  -(����  -(����  .����  .����  -(����      !    ,  0\����  0\����  18����  18����  0\����      !    ,����  h����  D��Ϥ  D��Ϥ  h����  h      !    ,����  h����  D����  D����  h����  h      !    ,��Ԯ  h��Ԯ  D��Պ  D��Պ  h��Ԯ  h      !    ,����  h����  D��ؾ  D��ؾ  h����  h      !    ,��ڔ  h��ڔ  D���p  D���p  h��ڔ  h      !    ,����  h����  D��ޤ  D��ޤ  h����  h      !    ,���z  h���z  D���V  D���V  h���z  h      !    ,���  h���  D���  D���  h���  h      !    ,���`  h���`  D���<  D���<  h���`  h      !    ,���  h���  D���p  D���p  h���  h      !    ,���F  h���F  D���"  D���"  h���F  h      !    ,���z  h���z  D���V  D���V  h���z  h      !    ,���,  h���,  D���  D���  h���,  h      !    ,���`  h���`  D���<  D���<  h���`  h      !    ,���  h���  D����  D����  h���  h      !    ,���F  h���F  D���"  D���"  h���F  h      !    ,����  h����  D����  D����  h����  h      !    ,������������������Ϥ������Ϥ������������      !    ,����������������������������������������      !    ,��Ԯ������Ԯ������Պ������Պ������Ԯ����      !    ,������������������ؾ������ؾ������������      !    ,��ڔ������ڔ�������p�������p������ڔ����      !    ,������������������ޤ������ޤ������������      !    ,���z�������z�������V�������V�������z����      !    ,�����������������������������������      !    ,���`�������`�������<�������<�������`����      !    ,�����������������p�������p�����������      !    ,���F�������F�������"�������"�������F����      !    ,���z�������z�������V�������V�������z����      !    ,���,�������,���������������������,����      !    ,���`�������`�������<�������<�������`����      !    ,�������������������������������������      !    ,���F�������F�������"�������"�������F����      !    ,����������������������������������������      !    ,������������   n��Ϥ   n��Ϥ������������      !    ,������������   n����   n����������������      !    ,��Ԯ������Ԯ   n��Պ   n��Պ������Ԯ����      !    ,������������   n��ؾ   n��ؾ������������      !    ,��ڔ������ڔ   n���p   n���p������ڔ����      !    ,������������   n��ޤ   n��ޤ������������      !    ,���z�������z   n���V   n���V�������z����      !    ,����������   n���   n��������������      !    ,���`�������`   n���<   n���<�������`����      !    ,����������   n���p   n���p�����������      !    ,���F�������F   n���"   n���"�������F����      !    ,���z�������z   n���V   n���V�������z����      !    ,���,�������,   n���   n����������,����      !    ,���`�������`   n���<   n���<�������`����      !    ,����������   n����   n���������������      !    ,���F�������F   n���"   n���"�������F����      !    ,������������   n����   n����������������      "    ,������������  H��ϩ  H��ϩ������������      "    ,������������  H����  H����������������      "    ,��ԩ������ԩ  H��Տ  H��Տ������ԩ����      "    ,������������  H����  H����������������      "    ,��ڏ������ڏ  H���u  H���u������ڏ����      "    ,������������  H��ީ  H��ީ������������      "    ,���u�������u  H���[  H���[�������u����      "    ,����������  H���  H��������������      "    ,���[�������[  H���A  H���A�������[����      "    ,����������  H���u  H���u�����������      "    ,���A�������A  H���'  H���'�������A����      "    ,���u�������u  H���[  H���[�������u����      "    ,���'�������'  H���  H����������'����      "    ,���[�������[  H���A  H���A�������[����      "    ,����������  H����  H���������������      "    ,���A�������A  H���'  H���'�������A����      "    ,������������  H����  H����������������      "    ,  '����  '  H    H  ����  '����      "    ,  �����  �  H  �  H  �����  �����      "    ,  ����    H  �  H  �����  ����      "    ,  	�����  	�  H  
�  H  
�����  	�����      "    ,  �����  �  H  �  H  �����  �����      "    ,  �����  �  H  �  H  �����  �����      "    ,  �����  �  H  �  H  �����  �����      "    ,  �����  �  H  q  H  q����  �����      "    ,  �����  �  H  �  H  �����  �����      "    ,  q����  q  H  W  H  W����  q����      "    ,  �����  �  H  �  H  �����  �����      "    ,  !W����  !W  H  "=  H  "=����  !W����      "    ,  $�����  $�  H  %q  H  %q����  $�����      "    ,  '=����  '=  H  (#  H  (#����  '=����      "    ,  *q����  *q  H  +W  H  +W����  *q����      "    ,  -#����  -#  H  .	  H  .	����  -#����      "    ,  0W����  0W  H  1=  H  1=����  0W����          ,�������$����  �  3,  �  3,���$�������$          ,���T  ����T  8���L  8���L  ����T  �          ,���:  ����:  8���2  8���2  ����:  �          ,���   ����   8���  8���  ����   �          ,���  ����  8����  8����  ����  �          ,����  �����  8����  8����  �����  �          ,����  �����  8����  8����  �����  �          ,���  ����  8����  8����  ����  �          ,����  �����  8����  8����  �����  �          ,����  �����  8  |  8  |  �����  �          ,  j  �  j  8  b  8  b  �  j  �          ,  
P  �  
P  8  H  8  H  �  
P  �          ,  6  �  6  8  .  8  .  �  6  �          ,    �    8    8    �    �          ,    �    8  �  8  �  �    �          ,  !�  �  !�  8  $�  8  $�  �  !�  �          ,  '�  �  '�  8  *�  8  *�  �  '�  �          ,  -�  �  -�  8  0�  8  0�  �  -�  �          ,�����������  �  2  �  2����������          ,���T�������T������L������L�������T����          ,���:�������:������2������2�������:����          ,��� ������� ������������������� ����          ,�����������������������������������          ,��������������������������������������          ,��������������������������������������          ,�����������������������������������          ,��������������������������������������          ,���������������  |���  |������������          ,  j����  j���  b���  b����  j����          ,  
P����  
P���  H���  H����  
P����          ,  6����  6���  .���  .����  6����          ,  ����  ���  ���  ����  ����          ,  ����  ���  ����  �����  ����          ,  !�����  !����  $����  $�����  !�����          ,  '�����  '����  *����  *�����  '�����          ,  -�����  -����  0����  0�����  -�����     �     �      nfet_03v3_FTUVLQ    �    ,���
������
  �  1�  �  1�������
���          ,��΂���W��΂  ����  �������W��΂���W          ,���h���W���h  ����  �������W���h���W          ,���N���W���N  �����  ��������W���N���W          ,���4���W���4  �����  ��������W���4���W          ,������W���  ����  �������W������W          ,��� ���W���   ����  �������W��� ���W          ,�������W����  �����  ��������W�������W          ,�������W����  ����h  ����h���W�������W          ,�������W����  �  N  �  N���W�������W          ,  ����W  �  �  4  �  4���W  ����W          ,  	~���W  	~  �    �  ���W  	~���W          ,  d���W  d  �     �   ���W  d���W          ,  J���W  J  �  �  �  ����W  J���W          ,  0���W  0  �  �  �  ����W  0���W          ,  !���W  !  �  %�  �  %����W  !���W          ,  &����W  &�  �  +�  �  +����W  &����W          ,  ,����W  ,�  �  1~  �  1~���W  ,����W           ,���T  I���T  ����L  ����L  I���T  I           ,���:  I���:  ����2  ����2  I���:  I           ,���   I���   ����  ����  I���   I           ,���  I���  �����  �����  I���  I           ,����  I����  �����  �����  I����  I           ,����  I����  �����  �����  I����  I           ,���  I���  �����  �����  I���  I           ,����  I����  �����  �����  I����  I           ,����  I����  �  |  �  |  I����  I           ,  j  I  j  �  b  �  b  I  j  I           ,  
P  I  
P  �  H  �  H  I  
P  I           ,  6  I  6  �  .  �  .  I  6  I           ,    I    �    �    I    I           ,    I    �  �  �  �  I    I           ,  !�  I  !�  �  $�  �  $�  I  !�  I           ,  '�  I  '�  �  *�  �  *�  I  '�  I           ,  -�  I  -�  �  0�  �  0�  I  -�  I           ,������������  I  2  I  2������������           ,���T���q���T�������L�������L���q���T���q           ,���:���q���:�������2�������2���q���:���q           ,��� ���q��� �����������������q��� ���q           ,������q����������������������q������q           ,�������q�����������������������q�������q           ,�������q�����������������������q�������q           ,������q����������������������q������q           ,�������q�����������������������q�������q           ,�������q��������  |����  |���q�������q           ,  j���q  j����  b����  b���q  j���q           ,  
P���q  
P����  H����  H���q  
P���q           ,  6���q  6����  .����  .���q  6���q           ,  ���q  ����  ����  ���q  ���q           ,  ���q  ����  �����  ����q  ���q           ,  !����q  !�����  $�����  $����q  !����q           ,  '����q  '�����  *�����  *����q  '����q           ,  -����q  -�����  0�����  0����q  -����q          ,���:���{���:  ����f  ����f���{���:���{          ,��� ���{���   ����L  ����L���{��� ���{          ,������{���  ����2  ����2���{������{          ,�������{����  ����  �������{�������{          ,�������{����  �����  ��������{�������{          ,������{���  �����  ��������{������{          ,������{���  �����  ��������{������{          ,�������{����  �����  ��������{�������{          ,���j���{���j  �   �  �   ����{���j���{          ,  P���{  P  �  |  �  |���{  P���{          ,  6���{  6  �  b  �  b���{  6���{          ,  ���{    �  H  �  H���{  ���{          ,  ���{    �  .  �  .���{  ���{          ,  ����{  �  �    �  ���{  ����{          ,  "����{  "�  �  #�  �  #����{  "����{          ,  (����{  (�  �  )�  �  )����{  (����{          ,  .����{  .�  �  /�  �  /����{  .����{      !    ,����   }����  Y��Ϥ  Y��Ϥ   }����   }      !    ,����   }����  Y����  Y����   }����   }      !    ,��Ԯ   }��Ԯ  Y��Պ  Y��Պ   }��Ԯ   }      !    ,����   }����  Y��ؾ  Y��ؾ   }����   }      !    ,��ڔ   }��ڔ  Y���p  Y���p   }��ڔ   }      !    ,����   }����  Y��ޤ  Y��ޤ   }����   }      !    ,���z   }���z  Y���V  Y���V   }���z   }      !    ,���   }���  Y���  Y���   }���   }      !    ,���`   }���`  Y���<  Y���<   }���`   }      !    ,���   }���  Y���p  Y���p   }���   }      !    ,���F   }���F  Y���"  Y���"   }���F   }      !    ,���z   }���z  Y���V  Y���V   }���z   }      !    ,���,   }���,  Y���  Y���   }���,   }      !    ,���`   }���`  Y���<  Y���<   }���`   }      !    ,���   }���  Y����  Y����   }���   }      !    ,���F   }���F  Y���"  Y���"   }���F   }      !    ,����   }����  Y����  Y����   }����   }      !    ,  ,   }  ,  Y    Y     }  ,   }      !    ,  �   }  �  Y  �  Y  �   }  �   }      !    ,     }    Y  �  Y  �   }     }      !    ,  	�   }  	�  Y  
�  Y  
�   }  	�   }      !    ,  �   }  �  Y  �  Y  �   }  �   }      !    ,  �   }  �  Y  �  Y  �   }  �   }      !    ,  �   }  �  Y  �  Y  �   }  �   }      !    ,  �   }  �  Y  l  Y  l   }  �   }      !    ,  �   }  �  Y  �  Y  �   }  �   }      !    ,  v   }  v  Y  R  Y  R   }  v   }      !    ,  �   }  �  Y  �  Y  �   }  �   }      !    ,  !\   }  !\  Y  "8  Y  "8   }  !\   }      !    ,  $�   }  $�  Y  %l  Y  %l   }  $�   }      !    ,  'B   }  'B  Y  (  Y  (   }  'B   }      !    ,  *v   }  *v  Y  +R  Y  +R   }  *v   }      !    ,  -(   }  -(  Y  .  Y  .   }  -(   }      !    ,  0\   }  0\  Y  18  Y  18   }  0\   }      !    ,������������������Ϥ������Ϥ������������      !    ,����������������������������������������      !    ,��Ԯ������Ԯ������Պ������Պ������Ԯ����      !    ,������������������ؾ������ؾ������������      !    ,��ڔ������ڔ�������p�������p������ڔ����      !    ,������������������ޤ������ޤ������������      !    ,���z�������z�������V�������V�������z����      !    ,�����������������������������������      !    ,���`�������`�������<�������<�������`����      !    ,�����������������p�������p�����������      !    ,���F�������F�������"�������"�������F����      !    ,���z�������z�������V�������V�������z����      !    ,���,�������,���������������������,����      !    ,���`�������`�������<�������<�������`����      !    ,�������������������������������������      !    ,���F�������F�������"�������"�������F����      !    ,����������������������������������������      !    ,  ,����  ,����  ����  ����  ,����      !    ,  �����  �����  �����  �����  �����      !    ,  ����  ����  �����  �����  ����      !    ,  	�����  	�����  
�����  
�����  	�����      !    ,  �����  �����  �����  �����  �����      !    ,  �����  �����  �����  �����  �����      !    ,  �����  �����  �����  �����  �����      !    ,  �����  �����  l����  l����  �����      !    ,  �����  �����  �����  �����  �����      !    ,  v����  v����  R����  R����  v����      !    ,  �����  �����  �����  �����  �����      !    ,  !\����  !\����  "8����  "8����  !\����      !    ,  $�����  $�����  %l����  %l����  $�����      !    ,  'B����  'B����  (����  (����  'B����      !    ,  *v����  *v����  +R����  +R����  *v����      !    ,  -(����  -(����  .����  .����  -(����      !    ,  0\����  0\����  18����  18����  0\����      "    ,�������a����  ���ϩ  ���ϩ���a�������a      "    ,�������a����  �����  ��������a�������a      "    ,��ԩ���a��ԩ  ���Տ  ���Տ���a��ԩ���a      "    ,�������a����  �����  ��������a�������a      "    ,��ڏ���a��ڏ  ����u  ����u���a��ڏ���a      "    ,�������a����  ���ީ  ���ީ���a�������a      "    ,���u���a���u  ����[  ����[���a���u���a      "    ,������a���  ����  �������a������a      "    ,���[���a���[  ����A  ����A���a���[���a      "    ,������a���  ����u  ����u���a������a      "    ,���A���a���A  ����'  ����'���a���A���a      "    ,���u���a���u  ����[  ����[���a���u���a      "    ,���'���a���'  ����  �������a���'���a      "    ,���[���a���[  ����A  ����A���a���[���a      "    ,������a���  �����  ��������a������a      "    ,���A���a���A  ����'  ����'���a���A���a      "    ,�������a����  �����  ��������a�������a      "    ,  '���a  '  �    �  ���a  '���a      "    ,  ����a  �  �  �  �  ����a  ����a      "    ,  ���a    �  �  �  ����a  ���a      "    ,  	����a  	�  �  
�  �  
����a  	����a      "    ,  ����a  �  �  �  �  ����a  ����a      "    ,  ����a  �  �  �  �  ����a  ����a      "    ,  ����a  �  �  �  �  ����a  ����a      "    ,  ����a  �  �  q  �  q���a  ����a      "    ,  ����a  �  �  �  �  ����a  ����a      "    ,  q���a  q  �  W  �  W���a  q���a      "    ,  ����a  �  �  �  �  ����a  ����a      "    ,  !W���a  !W  �  "=  �  "=���a  !W���a      "    ,  $����a  $�  �  %q  �  %q���a  $����a      "    ,  '=���a  '=  �  (#  �  (#���a  '=���a      "    ,  *q���a  *q  �  +W  �  +W���a  *q���a      "    ,  -#���a  -#  �  .	  �  .	���a  -#���a      "    ,  0W���a  0W  �  1=  �  1=���a  0W���a     �     �      (UNNAMED)  
  nfet_03v3_FTUVLQ �  B�         3"���� + = ,nfet_03v3_FTUVLQ_0   
  pfet_03v3_6DGS6C   3,  � + = ,pfet_03v3_6DGS6C_0      
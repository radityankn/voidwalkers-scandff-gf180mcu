magic
tech gf180mcuD
magscale 1 10
timestamp 1755194955
<< checkpaint >>
rect -2000 -4000 2005 1
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use inv  x1
timestamp 0
transform 1 0 2 0 1 -2000
box 0 0 1 1
use mux_tg  x2
timestamp 0
transform 1 0 0 0 1 -2000
box 0 0 1 1
use mux_tg  x3
timestamp 0
transform 1 0 1 0 1 -2000
box 0 0 1 1
use inv  x4
timestamp 0
transform 1 0 3 0 1 -2000
box 0 0 1 1
use inv  x5
timestamp 0
transform 1 0 4 0 1 -2000
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 1280 0 0 0 A
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 1280 0 0 0 B
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 1280 0 0 0 VSS
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 1280 0 0 0 S
port 5 nsew
<< end >>

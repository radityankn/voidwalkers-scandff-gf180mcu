** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrnq/sch/mux_2x1.sch
.subckt mux_2x1 A B VDD S VSS OUT
*.PININFO VDD:B OUT:O A:I B:I S:I VSS:B
x1 VDD S S_INV VSS inv
x2 VDD TG_OUT net1 VSS inv
x3 VDD net1 OUT VSS inv
x4 VDD S A TG_OUT S_INV VSS mux_tg
x5 VDD S_INV B TG_OUT S VSS mux_tg
.ends

* expanding   symbol:  cells/sdffrnq/sch/inv.sym # of pins=4
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrnq/sch/inv.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrnq/sch/inv.sch
.subckt inv VDD IN OUT VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
M2 OUT IN VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M1 OUT IN VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends


* expanding   symbol:  cells/sdffrnq/sch/mux_tg.sym # of pins=6
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrnq/sch/mux_tg.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrnq/sch/mux_tg.sch
.subckt mux_tg VDD P_GATE IN OUT N_GATE VSS
*.PININFO VDD:B VSS:B OUT:O IN:I P_GATE:I N_GATE:I
M1 IN N_GATE OUT VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M2 IN P_GATE OUT VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
.ends


magic
tech gf180mcuD
magscale 1 10
timestamp 1756235029
<< nmos >>
rect -440 -85 -380 85
rect -276 -85 -216 85
rect -112 -85 -52 85
rect 52 -85 112 85
rect 216 -85 276 85
rect 380 -85 440 85
<< ndiff >>
rect -528 72 -440 85
rect -528 -72 -515 72
rect -469 -72 -440 72
rect -528 -85 -440 -72
rect -380 -85 -276 85
rect -216 72 -112 85
rect -216 -72 -187 72
rect -141 -72 -112 72
rect -216 -85 -112 -72
rect -52 -85 52 85
rect 112 72 216 85
rect 112 -72 141 72
rect 187 -72 216 72
rect 112 -85 216 -72
rect 276 72 380 85
rect 276 -72 305 72
rect 351 -72 380 72
rect 276 -85 380 -72
rect 440 72 528 85
rect 440 -72 469 72
rect 515 -72 528 72
rect 440 -85 528 -72
<< ndiffc >>
rect -515 -72 -469 72
rect -187 -72 -141 72
rect 141 -72 187 72
rect 305 -72 351 72
rect 469 -72 515 72
<< polysilicon >>
rect -440 85 -380 129
rect -276 85 -216 129
rect -112 85 -52 129
rect 52 85 112 129
rect 216 85 276 129
rect 380 85 440 129
rect -440 -129 -380 -85
rect -276 -129 -216 -85
rect -112 -129 -52 -85
rect 52 -129 112 -85
rect 216 -129 276 -85
rect 380 -129 440 -85
<< metal1 >>
rect -515 72 -469 83
rect -515 -83 -469 -72
rect -187 72 -141 83
rect -187 -83 -141 -72
rect 141 72 187 83
rect 141 -83 187 -72
rect 305 72 351 83
rect 305 -83 351 -72
rect 469 72 515 83
rect 469 -83 515 -72
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.85 l 0.3 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>

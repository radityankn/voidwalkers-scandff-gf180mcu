* NGSPICE file created from mux_tg.ext - technology: gf180mcuD

.option scale=5n

.subckt mux_toplevel_postlayout VDD INPUT_1 VSS OUT INPUT_2 SELECTOR
X0 VDD.t1 a_n60_n80.t2 OUT.t0 VDD.t0 pfet_03v3 ad=22.1n pd=0.47m as=37.4n ps=0.9m w=340 l=60
X1 a_580_n190.t0 SELECTOR.t0 VDD.t3 VDD.t2 pfet_03v3 ad=37.4n pd=0.9m as=44.2n ps=0.94m w=340 l=60
X2 a_n60_n80.t0 a_130_n80.t4 VSS.t7 VSS.t6 nfet_03v3 ad=21.93n pd=0.598m as=11.05n ps=0.3m w=170 l=60
X3 a_130_n80.t3 SELECTOR.t1 INPUT_2.t1 VDD.t7 pfet_03v3 ad=22.1n pd=0.47m as=41.14n ps=0.922m w=340 l=60
X4 INPUT_1.t1 SELECTOR.t2 a_130_n80.t2 VSS.t5 nfet_03v3 ad=22.1n pd=0.6m as=11.05n ps=0.3m w=170 l=60
X5 a_580_n190.t1 SELECTOR.t3 VSS.t4 VSS.t3 nfet_03v3 ad=18.7n pd=0.56m as=22.1n ps=0.6m w=170 l=60
X6 VSS.t2 a_n60_n80.t3 OUT.t1 VSS.t1 nfet_03v3 ad=11.05n pd=0.3m as=18.7n ps=0.56m w=170 l=60
X7 a_130_n80.t1 a_580_n190.t2 INPUT_2.t0 VSS.t0 nfet_03v3 ad=11.05n pd=0.3m as=20.57n ps=0.582m w=170 l=60
X8 a_n60_n80.t1 a_130_n80.t5 VDD.t6 VDD.t5 pfet_03v3 ad=43.86n pd=0.938m as=22.1n ps=0.47m w=340 l=60
X9 INPUT_1.t0 a_580_n190.t3 a_130_n80.t0 VDD.t4 pfet_03v3 ad=44.2n pd=0.94m as=22.1n ps=0.47m w=340 l=60
C0 INPUT_1 VDD 0.06805f
C1 OUT VDD 0.20422f
C2 SELECTOR INPUT_2 0.01847f
C3 SELECTOR VDD 0.44409f
C4 INPUT_1 SELECTOR 0.05446f
C5 VDD INPUT_2 0.01849f
R0 a_n60_n80.n0 a_n60_n80.t2 43.9743
R1 a_n60_n80.n0 a_n60_n80.t3 19.0326
R2 a_n60_n80.t0 a_n60_n80.n1 8.88289
R3 a_n60_n80.n1 a_n60_n80.n0 8.221
R4 a_n60_n80.n1 a_n60_n80.t1 4.31776
R5 OUT OUT.t1 8.89575
R6 OUT OUT.t0 7.20731
R7 VDD.t4 VDD.t2 666.668
R8 VDD.t5 VDD.t7 625
R9 VDD.t7 VDD.t4 263.889
R10 VDD.t0 VDD.t5 263.889
R11 VDD.n2 VDD.t0 137.601
R12 VDD.n1 VDD.t3 5.06776
R13 VDD.n1 VDD.n0 2.8847
R14 VDD.n0 VDD.t6 1.33874
R15 VDD.n0 VDD.t1 1.33874
R16 VDD.n2 VDD.n1 0.13925
R17 VDD VDD.n2 0.1055
R18 SELECTOR.n1 SELECTOR.t1 57.1838
R19 SELECTOR.n0 SELECTOR.t0 41.3672
R20 SELECTOR.n2 SELECTOR.n1 31.7555
R21 SELECTOR.n0 SELECTOR.t3 16.4255
R22 SELECTOR.n1 SELECTOR.t2 16.4255
R23 SELECTOR SELECTOR.n2 8.06238
R24 SELECTOR.n2 SELECTOR.n0 3.2855
R25 a_580_n190.n0 a_580_n190.t2 94.8227
R26 a_580_n190.n0 a_580_n190.t3 75.1746
R27 a_580_n190.n1 a_580_n190.t1 9.06387
R28 a_580_n190.t0 a_580_n190.n1 4.11549
R29 a_580_n190.n1 a_580_n190.n0 0.4055
R30 a_130_n80.n1 a_130_n80.t4 31.0255
R31 a_130_n80.n1 a_130_n80.t5 26.7672
R32 a_130_n80.n2 a_130_n80.n1 25.0398
R33 a_130_n80.n2 a_130_n80.n0 7.00682
R34 a_130_n80.n3 a_130_n80.n2 2.55988
R35 a_130_n80.n0 a_130_n80.t2 2.40932
R36 a_130_n80.n0 a_130_n80.t1 2.40932
R37 a_130_n80.t0 a_130_n80.n3 1.33874
R38 a_130_n80.n3 a_130_n80.t3 1.33874
R39 VSS.t5 VSS.t3 2836.36
R40 VSS.t6 VSS.t0 2659.09
R41 VSS.t0 VSS.t5 1122.73
R42 VSS.t1 VSS.t6 1122.73
R43 VSS.n2 VSS.t1 719.491
R44 VSS.n1 VSS.t4 9.78718
R45 VSS.n1 VSS.n0 6.53501
R46 VSS.n0 VSS.t7 2.40932
R47 VSS.n0 VSS.t2 2.40932
R48 VSS.n2 VSS.n1 0.16175
R49 VSS VSS.n2 0.083
R50 INPUT_2 INPUT_2.t0 8.87218
R51 INPUT_2 INPUT_2.t1 6.95124
R52 INPUT_1 INPUT_1.t1 8.87218
R53 INPUT_1 INPUT_1.t0 4.40883
C6 INPUT_1 VSS 0.05754f
C7 INPUT_2 VSS 0.08253f
C8 OUT VSS 0.26279f
C9 SELECTOR VSS 0.74741f
C10 VDD VSS 4.16213f
.ends


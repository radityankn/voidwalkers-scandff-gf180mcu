VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER Via4
  TYPE CUT ;
END Via4

LAYER Via3
  TYPE CUT ;
END Via3

LAYER Via2
  TYPE CUT ;
END Via2

LAYER Via1
  TYPE CUT ;
END Via1

LAYER Nwell
  TYPE MASTERSLICE ;
END Nwell

LAYER Metal1
  TYPE ROUTING ;
END Metal1

LAYER Metal3
  TYPE ROUTING ;
END Metal3

LAYER Metal2
  TYPE ROUTING ;
END Metal2

LAYER Metal4
  TYPE ROUTING ;
END Metal4

LAYER Metal5
  TYPE ROUTING ;
END Metal5

LAYER Pwell
  TYPE MASTERSLICE ;
END Pwell

MACRO gf180mcu_voidwalkers_sc_sdffrnq_4
  CLASS BLOCK ;
  FOREIGN gf180mcu_voidwalkers_sc_sdffrnq_4 ;
  ORIGIN 8.450 -0.500 ;
  SIZE 27.650 BY 6.350 ;
  PIN VDD
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -8.450 3.250 19.200 6.850 ;
      LAYER Metal1 ;
        RECT -8.450 6.150 19.200 6.850 ;
        RECT -7.000 4.700 -6.645 6.150 ;
        RECT -3.100 4.950 -2.750 6.150 ;
        RECT 1.050 4.950 1.400 6.150 ;
        RECT 3.000 6.000 3.800 6.150 ;
        RECT 3.450 4.950 3.800 6.000 ;
        RECT -7.000 4.050 -6.650 4.700 ;
        RECT 7.300 4.050 7.650 6.150 ;
        RECT 10.900 4.050 11.250 6.150 ;
        RECT 17.400 4.050 17.750 6.150 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -8.450 2.700 19.200 3.250 ;
        RECT -8.450 2.600 9.800 2.700 ;
        RECT 10.450 2.600 10.750 2.700 ;
        RECT 11.400 2.600 11.700 2.700 ;
        RECT 12.100 2.600 19.200 2.700 ;
        RECT -8.450 0.500 19.200 2.600 ;
      LAYER Metal1 ;
        RECT -7.000 1.200 -6.645 2.470 ;
        RECT -4.850 1.200 -4.500 2.450 ;
        RECT -2.950 1.200 -2.600 2.350 ;
        RECT 1.050 1.200 1.400 2.100 ;
        RECT 3.450 1.200 3.800 2.450 ;
        RECT 5.400 1.200 5.750 2.450 ;
        RECT 7.300 1.200 7.650 2.450 ;
        RECT 10.900 1.200 11.250 2.450 ;
        RECT 17.400 1.200 17.750 2.450 ;
        RECT -8.450 0.500 19.200 1.200 ;
    END
  END VSS
  PIN A
    ANTENNADIFFAREA 1.542750 ;
    PORT
      LAYER Metal1 ;
        RECT 14.050 3.050 14.400 4.850 ;
        RECT 13.800 2.600 14.400 3.050 ;
        RECT 14.050 1.600 14.400 2.600 ;
    END
  END A
  PIN B
    ANTENNADIFFAREA 1.657500 ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 3.050 16.300 5.750 ;
        RECT 15.700 2.600 16.300 3.050 ;
        RECT 15.950 1.600 16.300 2.600 ;
    END
  END B
  PIN S
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 17.450 2.700 18.200 3.150 ;
    END
  END S
  PIN CLK
    ANTENNAGATEAREA 3.060000 ;
    PORT
      LAYER Metal1 ;
        RECT -1.700 4.100 0.350 4.700 ;
        RECT -1.700 3.300 -1.200 4.100 ;
        RECT 0.000 2.900 0.350 4.100 ;
        RECT 12.700 3.050 13.300 3.650 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 2.900 4.250 3.650 ;
    END
  END RN
  PIN Q
    ANTENNADIFFAREA 1.402500 ;
    PORT
      LAYER Metal1 ;
        RECT -7.950 3.750 -7.600 5.750 ;
        RECT -8.350 3.000 -7.600 3.750 ;
        RECT -7.950 1.600 -7.600 3.000 ;
    END
  END Q
  OBS
      LAYER Metal1 ;
        RECT -6.050 3.200 -5.700 5.750 ;
        RECT -5.450 5.100 -4.350 5.750 ;
        RECT -5.450 3.300 -5.050 5.100 ;
        RECT -7.350 2.700 -5.700 3.200 ;
        RECT -4.700 3.050 -4.350 5.100 ;
        RECT -2.500 4.950 -0.900 5.750 ;
        RECT 1.650 5.100 3.200 5.750 ;
        RECT 5.500 5.400 6.750 5.750 ;
        RECT -2.500 4.700 -2.200 4.950 ;
        RECT 1.650 4.700 2.000 5.100 ;
        RECT -3.650 4.400 -2.200 4.700 ;
        RECT 0.600 4.400 2.000 4.700 ;
        RECT -3.650 3.600 -3.100 4.400 ;
        RECT -3.650 3.300 -1.950 3.600 ;
        RECT -4.700 2.700 -2.450 3.050 ;
        RECT -6.050 1.600 -5.700 2.700 ;
        RECT -3.900 2.600 -2.450 2.700 ;
        RECT -3.900 1.600 -3.500 2.600 ;
        RECT -2.200 2.150 -1.950 3.300 ;
        RECT -0.750 2.650 -0.350 3.800 ;
        RECT 0.600 3.500 1.200 4.400 ;
        RECT 2.250 2.650 2.600 4.850 ;
        RECT 2.850 4.700 3.200 5.100 ;
        RECT 4.050 5.150 6.750 5.400 ;
        RECT 4.050 5.100 5.900 5.150 ;
        RECT 4.050 4.700 4.350 5.100 ;
        RECT 2.850 4.350 4.350 4.700 ;
        RECT 4.600 4.050 5.300 4.850 ;
        RECT 5.550 4.050 5.900 5.100 ;
        RECT 5.000 3.800 5.300 4.050 ;
        RECT 5.000 3.400 6.200 3.800 ;
        RECT 5.000 3.050 5.300 3.400 ;
        RECT -0.750 2.350 2.600 2.650 ;
        RECT -2.200 1.600 -0.900 2.150 ;
        RECT 2.000 1.600 2.600 2.350 ;
        RECT 4.600 2.700 5.300 3.050 ;
        RECT 6.450 3.150 6.750 5.150 ;
        RECT 7.900 5.150 9.350 5.750 ;
        RECT 7.900 3.800 8.250 5.150 ;
        RECT 7.000 3.400 8.250 3.800 ;
        RECT 6.450 2.700 8.300 3.150 ;
        RECT 4.600 1.600 4.950 2.700 ;
        RECT 6.450 2.450 6.750 2.700 ;
        RECT 6.350 1.600 6.750 2.450 ;
        RECT 9.000 1.600 9.350 5.150 ;
        RECT 11.500 5.100 15.350 5.750 ;
        RECT 11.500 3.800 11.850 5.100 ;
        RECT 10.450 3.500 11.850 3.800 ;
        RECT 12.100 3.150 12.450 4.850 ;
        RECT 9.600 2.700 12.450 3.150 ;
        RECT 12.100 2.450 12.450 2.700 ;
        RECT 11.850 1.600 12.450 2.450 ;
        RECT 15.000 1.600 15.350 5.100 ;
        RECT 16.750 3.800 17.150 5.900 ;
        RECT 18.350 4.050 18.900 5.750 ;
        RECT 18.600 3.800 18.900 4.050 ;
        RECT 16.750 3.400 18.900 3.800 ;
        RECT 16.750 1.450 17.150 3.400 ;
        RECT 18.600 2.450 18.900 3.400 ;
        RECT 18.350 1.600 18.900 2.450 ;
  END
END gf180mcu_voidwalkers_sc_sdffrnq_4
END LIBRARY


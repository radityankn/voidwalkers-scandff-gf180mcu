** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_toplevel.sch
**.subckt mux_toplevel vdd data vss out scan_data se_in
*.iopin vdd
*.opin out
*.ipin data
*.ipin scan_data
*.ipin se_in
*.iopin vdd
*.iopin vss
*.iopin vss
*.iopin vdd
*.iopin vss
x2 vdd net1 data net2 se_in vss mux_tg
x1 vdd se_in net1 vss mux_inverter
x3 vdd se_in scan_data net2 net1 vss mux_tg
x4 vdd net2 net3 vss mux_inverter
x5 vdd net3 out vss mux_inverter
**.ends

* expanding   symbol:  voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_tg.sym # of pins=6
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_tg.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_tg.sch
.subckt mux_tg VDD P_GATE IN OUT N_GATE VSS
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin IN
*.ipin P_GATE
*.ipin N_GATE
XM1 IN N_GATE OUT VSS nfet_03v3 L=0.3u W=0.85u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 IN P_GATE OUT VDD pfet_03v3 L=0.3u W=1.7u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_inverter.sym # of pins=4
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_inverter.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_inverter.sch
.subckt mux_inverter vdd in out_inv gnd
*.iopin vdd
*.iopin gnd
*.opin out_inv
*.ipin in
XM1 out_inv in gnd gnd nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 out_inv in vdd vdd pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.end

magic
tech gf180mcuD
magscale 1 10
timestamp 1756235029
<< nwell >>
rect 0 585 3038 1270
<< psubdiff >>
rect 49 121 194 140
rect 49 72 89 121
rect 155 72 194 121
rect 2020 117 2165 139
rect 49 48 194 72
rect 2020 68 2062 117
rect 2128 68 2165 117
rect 2020 47 2165 68
rect 2322 117 2467 139
rect 2322 68 2364 117
rect 2430 68 2467 117
rect 2322 47 2467 68
rect 2588 118 2733 140
rect 2588 69 2628 118
rect 2694 69 2733 118
rect 2588 48 2733 69
rect 2891 121 3036 140
rect 2891 72 2930 121
rect 2996 72 3036 121
rect 2891 48 3036 72
<< nsubdiff >>
rect 58 1199 203 1222
rect 58 1150 98 1199
rect 164 1150 203 1199
rect 1940 1198 2085 1222
rect 58 1130 203 1150
rect 1940 1149 1978 1198
rect 2044 1149 2085 1198
rect 1940 1130 2085 1149
rect 2223 1194 2368 1221
rect 2223 1145 2264 1194
rect 2330 1145 2368 1194
rect 2223 1129 2368 1145
rect 2502 1197 2647 1222
rect 2502 1148 2543 1197
rect 2609 1148 2647 1197
rect 2502 1130 2647 1148
rect 2777 1196 2922 1219
rect 2777 1149 2821 1196
rect 2887 1149 2922 1196
rect 2777 1129 2922 1149
<< psubdiffcont >>
rect 89 72 155 121
rect 2062 68 2128 117
rect 2364 68 2430 117
rect 2628 69 2694 118
rect 2930 72 2996 121
<< nsubdiffcont >>
rect 98 1150 164 1199
rect 1978 1149 2044 1198
rect 2264 1145 2330 1194
rect 2543 1148 2609 1197
rect 2821 1149 2887 1196
<< polysilicon >>
rect 534 1158 1511 1218
rect 736 51 1578 111
<< metal1 >>
rect 1298 611 1619 671
<< metal2 >>
rect 1269 834 2266 894
rect 1269 534 1329 834
rect 2326 477 2427 537
rect 533 282 1685 342
use dff  dff_0
timestamp 1756208311
transform 1 0 0 0 1 423
box 0 -423 1551 847
use dff_1  dff_1_0
timestamp 1756235029
transform 1 0 1112 0 1 423
box 236 -423 1932 847
<< labels >>
flabel space 304 516 309 518 0 FreeSans 240 0 0 0 CLK
port 0 nsew
flabel nwell 463 636 468 638 0 FreeSans 240 0 0 0 D
port 1 nsew
flabel nwell 47 1194 48 1195 0 FreeSans 240 0 0 0 VDD
port 2 nsew
flabel psubdiff 52 57 52 57 0 FreeSans 240 0 0 0 VSS
port 3 nsew
flabel space 1300 510 1300 510 0 FreeSans 240 0 0 0 R
port 4 nsew
flabel space 2996 546 2996 546 0 FreeSans 240 0 0 0 Q
port 5 nsew
<< end >>

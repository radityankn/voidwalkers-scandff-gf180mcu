  X � 	   & )� 	   & ) sdffrnq  >A�7KƧ�9D�/��ZT � 	   & )� 	   & ) mux_as_component        ,  r  �  r  �  ~  �  ~  �  r  �      �    ,  r���  r  �  ~  �  ~���  r���          ,  �  �  �  �  �  �  �  �  �  �          ,  �  �  �  �  �  �  �  �  �  �          ,  ����j  �  �  �  �  ����j  ����j          ,  ����j  �  �  �  �  ����j  ����j           ,  
n  \  
n  �    �    \  
n  \           ,  �  \  �  �  |  �  |  \  �  \           ,  W����  W  \  `  \  `����  W����           ,  @����  @  \  \  \  \����  @����           ,  
n����  
n����  ����  ����  
n����           ,  �����  �����  |����  |����  �����          ,  
n  @  
n  �    �    @  
n  @          ,  �  @  �  �  |  �  |  @  �  @          ,  W  \  W  @  `  @  `  \  W  \          ,  @  \  @  @  \  @  \  \  @  \          ,  
n    
n  \    \      
n            ,  �    �  \  |  \  |    �            ,  
  �  
  �  |  �  |  �  
  �          ,  T    T  �  �  �  �    T            ,  
    
  �  6  �  6    
            ,  �  �  �  �  |  �  |  �  �  �          ,  T  �  T    6    6  �  T  �          ,  
  �  
  �  6  �  6  �  
  �          ,  j  �  j  �  �  �  �  �  j  �          ,  
  �  
  �  �  �  �  �  
  �          ,  T���v  T  �  �  �  ����v  T���v          ,  
���p  
  �  6  �  6���p  
���p          ,  ����v  �  ^  |  ^  |���v  ����v          ,  j���p  j  �  �  �  ����p  j���p          ,  T���J  T���v  |���v  |���J  T���J      !    ,  F  �  F  �  "  �  "  �  F  �      !    ,  W  �  W  ~  3  ~  3  �  W  �      !    ,    �    ~  �  ~  �  �    �      !    ,  �  �  �  ~  �  ~  �  �  �  �      !    ,  m  �  m  ~  I  ~  I  �  m  �      !    ,  	�  
  	�  
�  
}  
�  
}  
  	�  
      !    ,  W  
  W  
�  3  
�  3  
  W  
      !    ,    
    
�  �  
�  �  
    
      !    ,  �  
  �  
�  �  
�  �  
  �  
      !    ,  m  
  m  
�  I  
�  I  
  m  
      !    ,  �  B  �    �    �  B  �  B      !    ,  	�   �  	�  �  
}  �  
}   �  	�   �      !    ,  W   �  W  �  3  �  3   �  W   �      !    ,     �    �  �  �  �   �     �      !    ,  �   �  �  �  �  �  �   �  �   �      !    ,  m   �  m  �  I  �  I   �  m   �      !    ,  F���t  F   P  "   P  "���t  F���t      "    ,  r  �  r  �  ~  �  ~  �  r  �      "    ,  r    r  �  t  �  t    r        "    ,  	`    	`    
�    
�    	`        "    ,  f  R  f    
�    
�  R  f  R      "    ,  	`���j  	`  R  
�  R  
����j  	`���j      "    ,  ���j      t    t���j  ���j      "    ,  �    �  �  *  �  *    �        "    ,  �  R  �    *    *  R  �  R      "    ,  ����j  �  R  *  R  *���j  ����j      "    ,  �    �  �  |  �  |    �        "    ,  v  �  v  �  �  �  �  �  v  �      "    ,  ,  �  ,  �  R  �  R  �  ,  �      "    ,  &    &  �  R  �  R    &        "    ,  �  r  �    R    R  r  �  r      "    ,  ����p  �  r  |  r  |���p  ����p      "    ,  �  �  �  x  �  x  �  �  �  �      "    ,  &  �  &  r  R  r  R  �  &  �      "    ,  v���v  v  �  �  �  ����v  v���v      "    ,  ,���j  ,  �  R  �  R���j  ,���j      "    ,  r���  r���v  ~���v  ~���  r���     � 	   & )� 	   & ) sdffrnq  
  mux_as_component   -�  � + = ,mux_as_component_0          ,����  �����  �  3�  �  3�  �����  �      �    ,����  
�����  �  3�  �  3�  
�����  
�      �    ,����  
(����  
�  &H  
�  &H  
(����  
(      �    ,  (�  
(  (�  
�  )�  
�  )�  
(  (�  
(      �    ,  ,�  
(  ,�  
�  -�  
�  -�  
(  ,�  
(      �    ,  /D  
(  /D  
�  3�  
�  3�  
(  /D  
(      �    ,����  �����  
(  3�  
(  3�  �����  �          ,����  j����  ,����  ,����  j����  j          ,  �  p  �  2  t  2  t  p  �  p          ,  .J  j  .J  ,  2�  ,  2�  j  .J  j          ,����  �����  v���M  v���M  �����  �          ,���r  ����r  v  
�  v  
�  ����r  �          ,  H  �  H  D  �  D  �  �  H  �          ,  |  �  |  v  18  v  18  �  |  �          ,����  @����  	����M  	����M  @����  @          ,����  @����  	�  
�  	�  
�  @����  @          ,  H  @  H  	�  �  	�  �  @  H  @          ,  �  @  �  	�  18  	�  18  @  �  @          ,����  �����  L���  L���  �����  �          ,����  �����  L���  L���  �����  �          ,����  �����  L���j  L���j  �����  �          ,  .J  �  .J  L  2�  L  2�  �  .J  �           ,���   t���   ����  ����  t���   t           ,    t    �    �    t    t           ,  -�  t  -�  �  3�  �  3�  t  -�  t           ,���  V���  t����  t����  V���  V           ,  �  \  �  t  �  t  �  \  �  \           ,  .6  V  .6  t  3�  t  3�  V  .6  V           ,  1�  �  1�  V  3�  V  3�  �  1�  �           ,���   
2���   
x���  
x���  
2���   
2           ,���  
2���  
x���n  
x���n  
2���  
2           ,���L  
2���L  
x     
x     
2���L  
2           ,  �  
2  �  
x  �  
x  �  
2  �  
2           ,  &  
2  &  
x  .�  
x  .�  
2  &  
2           ,���   ����   
2  1�  
2  1�  ����   �           ,���   Z���   ����  ����  Z���   Z           ,���  Z���  ����n  ����n  Z���  Z           ,���L  Z���L  �     �     Z���L  Z           ,  �  Z  �  �  �  �  �  Z  �  Z           ,  &  Z  &  �  .�  �  .�  Z  &  Z          ,���   ���   \���  \���  ���             ,���  ���  \����  \����  ���            ,����  ����  \���$  \���$  ����            ,  r    r  \     \       r            ,���   2���   ����  ����  2���   2          ,����  �����    ^    ^  �����  �          ,  �  �  �  *  �  *  �  �  �  �          ,  �    �  \  .�  \  .�    �            ,  �  �  �    1�    1�  �  �  �          ,����  2����  �  1�  �  1�  2����  2          ,���   ����   2���  2���  ����   �          ,���  ����  2����  2����  ����  �          ,����  �����  2���$  2���$  �����  �          ,  r  �  r  2     2     �  r  �          ,  �     �  2  (  2  (     �             ,  �  �  �     �     �  �  �  �          ,  �  �  �  2  .�  2  .�  �  �  �          ,��߲  v��߲  `���  `���  v��߲  v          ,���  v���  `���  `���  v���  v          ,����  v����  `���~  `���~  v����  v          ,  .6  v  .6  `  3  `  3  v  .6  v          ,���  ����  ^  �  ^  �  ����  �          ,����  �����  p���  p���  �����  �          ,���  ����  p����  p����  ����  �          ,���  <���  �����  �����  <���  <          ,���  ����  ����  ����  ����  �          ,���  ����  <����  <����  ����  �          ,���  <���  p����  p����  <���  <          ,���n  <���n  p����  p����  <���n  <          ,���  ���  <����  <����  ���            ,���  ���  <����  <����  ���            ,���\  <���\  p����  p����  <���\  <          ,����  
�����  ����  ����  
�����  
�          ,����  F����  
����  
����  F����  F          ,���  F���  �����  �����  F���  F          ,���  F���  ����.  ����.  F���  F          ,���  T���  ����  ����  T���  T          ,���  ����  ���n  ���n  ����  �          ,���\  ����\  <���P  <���P  ����\  �          ,���  ����  p���>  p���>  ����  �          ,  X  <  X  p  �  p  �  <  X  <          ,����  N����  �����  �����  N����  N          ,���  
(���  T����  T����  
(���  
(          ,���  
(���  �����  �����  
(���  
(          ,���  T���  N���>  N���>  T���  T          ,���  F���  
(����  
(����  F���  F          ,���n  F���n  
(����  
(����  F���n  F          ,���\  
(���\  T���>  T���>  
(���\  
(          ,����  
�����  �  ^  �  ^  
�����  
�          ,���\  F���\  
(����  
(����  F���\  F          ,   2  L   2  
�  ^  
�  ^  L   2  L          ,  X  H  X  <  �  <  �  H  X  H          ,  X  F  X  H  �  H  �  F  X  F          ,    L    p  :  p  :  L    L          ,  n  B  n  p  �  p  �  B  n  B          ,  �  <  �  �  �  �  �  <  �  <          ,  %  j  %  �  -�  �  -�  j  %  j          ,  �  T  �  B  �  B  �  T  �  T          ,  �  �  �  <  �  <  �  �  �  �          ,  �  <  �  p  �  p  �  <  �  <          ,  �    �  <  ~  <  ~    �            ,  n  F  n  T  �  T  �  F  n  F          ,    F    �  8  �  8  F    F          ,  �  F  �    �    �  F  �  F          ,  x  �  x  p  �  p  �  �  x  �          ,  !f  �  !f  p  "�  p  "�  �  !f  �          ,  %  �  %  j  &H  j  &H  �  %  �          ,  (�  <  (�  p  )�  p  )�  <  (�  <          ,  !f  �  !f  �  &H  �  &H  �  !f  �          ,  x  
�  x  �   l  �   l  
�  x  
�          ,  %  N  %  �  &H  �  &H  N  %  N          ,  (�  H  (�  <  +*  <  +*  H  (�  H          ,  ,�  �  ,�  j  -�  j  -�  �  ,�  �          ,  1�  �  1�  B  3�  B  3�  �  1�  �          ,  %  
�  %  N  't  N  't  
�  %  
�          ,  x  F  x  
�  �  
�  �  F  x  F          ,  !f  L  !f  
�  "�  
�  "�  L  !f  L          ,  %  F  %  
�  &H  
�  &H  F  %  F          ,  (�  F  (�  H  )�  H  )�  F  (�  F          ,  ,�  �  ,�  �  3�  �  3�  �  ,�  �          ,  ,�  L  ,�  �  -�  �  -�  L  ,�  L          ,  1�  �  1�  �  3�  �  3�  �  1�  �          ,   2      2  L  -�  L  -�      2         !    ,����  �����  ����  ����  �����  �      !    ,  /I  �  /I  �  0%  �  0%  �  /I  �      !    ,  1  �  1  �  1�  �  1�  �  1  �      !    ,  �  �  �  �  �  �  �  �  �  �      !    ,���3  x���3  T���  T���  x���3  x      !    ,����  x����  T����  T����  x����  x      !    ,���  x���  T���{  T���{  x���  x      !    ,����  x����  T����  T����  x����  x      !    ,���%  x���%  T���  T���  x���%  x      !    ,���-  x���-  T���	  T���	  x���-  x      !    ,  [  x  [  T  7  T  7  x  [  x      !    ,  �  F  �  "  �  "  �  F  �  F      !    ,  �  x  �  T  �  T  �  x  �  x      !    ,  �  x  �  T  �  T  �  x  �  x      !    ,  #i  x  #i  T  $E  T  $E  x  #i  x      !    ,  *�  x  *�  T  +�  T  +�  x  *�  x      !    ,����  �����  �����  �����  �����  �      !    ,���  ����  ����{  ����{  ����  �      !    ,����  �����  �����  �����  �����  �      !    ,  	  �  	  �  	�  �  	�  �  	  �      !    ,  9  �  9  �    �    �  9  �      !    ,  �  �  �  �  �  �  �  �  �  �      !    ,  �  �  �  �  �  �  �  �  �  �      !    ,  #i  �  #i  �  $E  �  $E  �  #i  �      !    ,  *�  �  *�  �  +�  �  +�  �  *�  �      !    ,  /�  �  /�  �  0a  �  0a  �  /�  �      !    ,���  p���  L����  L����  p���  p      !    ,���c  ����c  ����?  ����?  ����c  �      !    ,����  �����  ~����  ~����  �����  �      !    ,���:  %���:  ���  ���  %���:  %      !    ,     W     3   �  3   �  W     W      !    ,    �    �  �  �  �  �    �      !    ,  �  �  �  ~  a  ~  a  �  �  �      !    ,  �  �  �  �  �  �  �  �  �  �      !    ,  )�  �  )�  �  *l  �  *l  �  )�  �      !    ,  �  ]  �  9  �  9  �  ]  �  ]      !    ,  2Z  �  2Z  �  36  �  36  �  2Z  �      !    ,����  ����  ����  ����  ����        !    ,����  
�����  w���_  w���_  
�����  
�      !    ,    1      �    �  1    1      !    ,  %�  
�  %�  �  &�  �  &�  
�  %�  
�      !    ,���3  {���3  W���  W���  {���3  {      !    ,����  {����  W����  W����  {����  {      !    ,���  {���  W���{  W���{  {���  {      !    ,���O  {���O  W���+  W���+  {���O  {      !    ,���  {���  W����  W����  {���  {      !    ,����  I����  %����  %����  I����  I      !    ,���-  ���-  ����	  ����	  ���-        !    ,  [  �  [  �  7  �  7  �  [  �      !    ,    {    W  �  W  �  {    {      !    ,  �  {  �  W  �  W  �  {  �  {      !    ,  9  {  9  W    W    {  9  {      !    ,  Y  {  Y  W  5  W  5  {  Y  {      !    ,    {    W  �  W  �  {    {      !    ,  �  {  �  W  �  W  �  {  �  {      !    ,  #i  {  #i  W  $E  W  $E  {  #i  {      !    ,  *�  {  *�  W  +�  W  +�  {  *�  {      !    ,  .�  {  .�  W  /g  W  /g  {  .�  {      !    ,���  ����  ����  ����  ����  �      !    ,����  �����  ����  ����  �����  �      !    ,���  ����  ����  ����  ����  �      !    ,����  �����  �����  �����  �����  �      !    ,����  �����  ����k  ����k  �����  �      !    ,  /I  �  /I  �  0%  �  0%  �  /I  �      !    ,  1  �  1  �  1�  �  1�  �  1  �      "    ,����  j����  �  3�  �  3�  j����  j      "    ,����  �����  v���P  v���P  �����  �      "    ,���  \���  j���  j���  \���  \      "    ,���  ����  \���  \���  ����  �      "    ,���b  ����b  ����P  ����P  ����b  �      "    ,���^  ����^  v���  v���  ����^  �      "    ,���  ����  v���  v���  ����  �      "    ,���  ����  ����F  ����F  ����  �      "    ,����  @����  ����P  ����P  @����  @      "    ,���J  
����J  ����  ����  
����J  
�      "    ,���  ����  ����  ����  ����  �      "    ,����  V����  j���B  j���B  V����  V      "    ,���<  V���<  v���|  v���|  V���<  V      "    ,    V    j  x  j  x  V    V      "    ,  �  p  �  j  �  j  �  p  �  p      "    ,  r  �  r  v  �  v  �  �  r  �      "    ,���<  \���<  V���h  V���h  \���<  \      "    ,  r  \  r  �  �  �  �  \  r  \      "    ,���  0���  \���h  \���h  0���  0      "    ,���  ���  0����  0����  ���        "    ,���\  ���\  \  ^  \  ^  ���\        "    ,���  ����  ���b  ���b  ����  �      "    ,���\  ����\  ���P  ���P  ����\  �      "    ,���  
����  ����n  ����n  
����  
�      "    ,���  L���  	����  	����  L���  L      "    ,���^  @���^  
����  
����  @���^  @      "    ,����  
(����  
����n  
����n  
(����  
(      "    ,���  L���  	����l  	����l  L���  L      "    ,����  @����  
(���T  
(���T  @����  @      "    ,���z  L���z  	.����  	.����  L���z  L      "    ,���h  f���h  ����b  ����b  f���h  f      "    ,���  
Z���  �����  �����  
Z���  
Z      "    ,      T        ^    ^  T      T      "    ,  X  0  X  \  �  \  �  0  X  0      "    ,  X  �  X  0  �  0  �  �  X  �      "    ,  �  
Z  �  �  
(  �  
(  
Z  �  
Z      "    ,  "  \  "  �  �  �  �  \  "  \      "    ,  z  V  z  p  �  p  �  V  z  V      "    ,  |    |  v  ^  v  ^    |        "    ,  �    �    ^    ^    �        "    ,  �  �  �          �  �  �      "    ,  �  \  �  �  �  �  �  \  �  \      "    ,  "  �  "  \  �  \  �  �  "  �      "    ,  �  �  �  �  �  �  �  �  �  �      "    ,  �  �  �  �    �    �  �  �      "    ,  �  �  �  �  �  �  �  �  �  �      "    ,  �  T  �  B  �  B  �  T  �  T      "    ,  �  H  �  �  8  �  8  H  �  H      "    ,  �  �  �  H  �  H  �  �  �  �      "    ,���  	.���  
Z  
(  
Z  
(  	.���  	.      "    ,  �  
�  �  �  �  �  �  
�  �  
�      "    ,  2  N  2    ^    ^  N  2  N      "    ,  �  �  �  j  �  j  �  �  �  �      "    ,  �    �  v  $�  v  $�    �        "    ,  �  �  �     :     :  �  �  �      "    ,  X  H  X  �   :  �   :  H  X  H      "    ,  2  
�  2  N   l  N   l  
�  2  
�      "    ,���h  @���h  f���|  f���|  @���h  @      "    ,    L    4  x  4  x  L    L      "    ,  �  @  �  	.  
(  	.  
(  @  �  @      "    ,  z  L  z  	�  �  	�  �  L  z  L      "    ,  �  @  �  
�  V  
�  V  @  �  @      "    ,  2  	�  2  
�  ^  
�  ^  	�  2  	�      "    ,    L    	�  v  	�  v  L    L      "    ,  �  @  �  	�  ^  	�  ^  @  �  @      "    ,  �  L  �  	�  �  	�  �  L  �  L      "    ,  #(  @  #(    $�    $�  @  #(  @      "    ,  *�  �  *�  j  +�  j  +�  �  *�  �      "    ,  ,�  �  ,�  v  3�  v  3�  �  ,�  �      "    ,  ,�  �  ,�  �  .J  �  .J  �  ,�  �      "    ,  (�  �  (�  �  .J  �  .J  �  (�  �      "    ,  /D  N  /D  �  0�  �  0�  N  /D  N      "    ,  %�  
�  %�  N  0�  N  0�  
�  %�  
�      "    ,  1�  �  1�  B  3�  B  3�  �  1�  �      "    ,  /D  	�  /D  
�  0�  
�  0�  	�  /D  	�      "    ,  *�  L  *�  	�  +�  	�  +�  L  *�  L      "    ,  .J  @  .J  	�  0�  	�  0�  @  .J  @      "    ,����  �����  L  3�  L  3�  �����  �      "  
 ,����  j����  �  K   �  K   j����  j      "  
 ,����  �����  L  K   L  K   �����  �      "  
 ,  5�  
(  5�  �  8@  �  8@  
(  5�  
(      "  
 ,  =T  
(  =T  �  ?�  �  ?�  
(  =T  
(      "  
 ,  D*  
�  D*  N  G  N  G  
�  D*  
�      "  
 ,  1�  �  1�  B  3�  B  3�  �  1�  �      "  
 ,  �  T  �  B  �  B  �  T  �  T      "  
 ,���b  ����b  ����P  ����P  ����b  �      "  
      @L������   �  � VDD       "  
      @L������   �    VSS       "  
      @L������   7  	 A       "  
      @L������   >�  	 B       "  
      @L������   E�  m S       "  
      @L������   2�   CLK       "  
      @L������   #  � RN      "  
      @L������ ����  / Q       
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrnq/sch/d_flip_flop_r.sch
.subckt d_flip_flop_r VDD VSS Q D CLK RN
*.PININFO D:I VDD:I VSS:I Q:O CLK:I RN:I
M1 net1 D VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M2 PROBE[0] CLK_INV net2 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M3 PROBE[0] CLK net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M4 net2 D VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M5 CLK_INV CLK VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M8 CLK_INV CLK VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M13 net3 PROBE[1] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M14 PROBE[0] CLK net4 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M15 PROBE[0] CLK_INV net3 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M16 net4 PROBE[1] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M9 net5 PROBE[1] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M10 PROBE[2] CLK net6 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M11 PROBE[2] CLK_INV net5 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M12 net6 PROBE[1] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M19 net7 PROBE[3] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M20 PROBE[2] CLK_INV net8 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M21 PROBE[2] CLK net7 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M22 net8 PROBE[3] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M23 QN PROBE[3] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M24 QN PROBE[3] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M25 Q QN VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M26 Q QN VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M6 net9 PROBE[0] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M27 PROBE[1] R net9 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M28 PROBE[1] PROBE[0] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M17 net10 PROBE[2] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M29 PROBE[3] R net10 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M30 PROBE[3] PROBE[2] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M7 PROBE[1] R VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M18 PROBE[3] R VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M31 R RN VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M32 R RN VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends

magic
tech gf180mcuD
magscale 1 10
timestamp 1756652194
<< nwell >>
rect -260 300 450 1020
<< pwell >>
rect -260 -250 450 300
<< nmos >>
rect -60 -30 0 140
rect 130 -30 190 140
<< pmos >>
rect -60 460 0 800
rect 130 460 190 800
<< ndiff >>
rect -170 120 -60 140
rect -170 -10 -150 120
rect -100 -10 -60 120
rect -170 -30 -60 -10
rect 0 120 130 140
rect 0 -10 40 120
rect 90 -10 130 120
rect 0 -30 130 -10
rect 190 120 319 140
rect 190 -10 230 120
rect 280 -10 319 120
rect 190 -30 319 -10
<< pdiff >>
rect -170 780 -60 800
rect -170 660 -150 780
rect -100 660 -60 780
rect -170 460 -60 660
rect 0 780 130 800
rect 0 660 40 780
rect 90 660 130 780
rect 0 600 130 660
rect 0 480 40 600
rect 90 480 130 600
rect 0 460 130 480
rect 190 780 319 800
rect 190 660 230 780
rect 280 660 319 780
rect 190 600 319 660
rect 190 480 230 600
rect 280 480 319 600
rect 190 460 319 480
<< ndiffc >>
rect -150 -10 -100 120
rect 40 -10 90 120
rect 230 -10 280 120
<< pdiffc >>
rect -150 660 -100 780
rect 40 660 90 780
rect 40 480 90 600
rect 230 660 280 780
rect 230 480 280 600
<< psubdiff >>
rect -220 -150 -80 -130
rect -220 -200 -200 -150
rect -100 -200 -80 -150
rect -220 -220 -80 -200
<< nsubdiff >>
rect -170 970 -70 990
rect -170 920 -150 970
rect -90 920 -70 970
rect -170 900 -70 920
<< psubdiffcont >>
rect -200 -200 -100 -150
<< nsubdiffcont >>
rect -150 920 -90 970
<< polysilicon >>
rect -60 800 0 850
rect 130 800 190 850
rect -60 290 0 460
rect 130 410 190 460
rect 130 390 440 410
rect 130 330 340 390
rect 420 330 440 390
rect 130 310 440 330
rect -60 270 80 290
rect -60 210 -40 270
rect 60 210 80 270
rect -60 190 80 210
rect -60 140 0 190
rect 130 140 190 310
rect -60 -80 0 -30
rect 130 -80 190 -30
<< polycontact >>
rect 340 330 420 390
rect -40 210 60 270
<< metal1 >>
rect -260 970 450 1020
rect -260 920 -150 970
rect -90 920 450 970
rect -260 900 450 920
rect -160 780 -90 800
rect -160 660 -150 780
rect -100 660 -90 780
rect -160 120 -90 660
rect 30 780 101 900
rect 30 660 40 780
rect 90 660 101 780
rect 30 600 101 660
rect 30 480 40 600
rect 90 590 101 600
rect 220 780 290 800
rect 220 660 230 780
rect 280 660 290 780
rect 220 600 290 660
rect 90 480 100 590
rect 30 460 100 480
rect 220 480 230 600
rect 280 480 290 600
rect 220 290 290 480
rect 340 670 450 800
rect 340 390 420 670
rect 340 310 420 330
rect -40 270 290 290
rect 60 210 290 270
rect -40 190 290 210
rect -160 -10 -150 120
rect -100 -10 -90 120
rect -160 -30 -90 -10
rect 30 120 101 144
rect 30 -10 40 120
rect 90 -10 101 120
rect 30 -130 101 -10
rect 220 120 290 190
rect 220 -10 230 120
rect 280 -10 290 120
rect 220 -30 290 -10
rect -260 -150 450 -130
rect -260 -200 -200 -150
rect -100 -200 450 -150
rect -260 -250 450 -200
<< end >>

** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_toplevel.sch
.subckt mux_toplevel vdd INPUT_1 vss out INPUT_2 SELECTOR
*.PININFO vdd:B out:O INPUT_1:I INPUT_2:I SELECTOR:I vdd:B vss:B vss:B vdd:B vss:B
x2 vdd net1 INPUT_1 net2 SELECTOR vss mux_tg
x1 vdd SELECTOR net1 vss mux_inverter
x3 vdd SELECTOR INPUT_2 net2 net1 vss mux_tg
x4 vdd net2 net3 vss mux_inverter
x5 vdd net3 out vss mux_inverter
.ends

* expanding   symbol:  voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_tg.sym # of pins=6
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_tg.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_tg.sch
.subckt mux_tg VDD P_GATE IN OUT N_GATE VSS
*.PININFO VDD:B VSS:B OUT:O IN:I P_GATE:I N_GATE:I
XM1 IN N_GATE OUT VSS nfet_03v3 L=0.3u W=0.85u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 IN P_GATE OUT VDD pfet_03v3 L=0.3u W=1.7u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_inverter.sym # of pins=4
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_inverter.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/libs/mux2x1_transmission_gate/mux_inverter.sch
.subckt mux_inverter vdd in out_inv gnd
*.PININFO vdd:B gnd:B out_inv:O in:I
XM1 out_inv in gnd gnd nfet_03v3 L=0.3u W=0.85u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 out_inv in vdd vdd pfet_03v3 L=0.3u W=1.7u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends


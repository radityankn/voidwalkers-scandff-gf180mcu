** sch_path: /foss/designs/libs/core_analog/unit_pmos/unit_pmos.sch
**.subckt unit_pmos drain sub gate source
*.iopin drain
*.iopin source
*.iopin sub
*.iopin gate
XM3 drain gate source sub pfet_03v3 L=0.5u W=8u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m={M}
**** begin user architecture code

.param M=1

**** end user architecture code
**.ends
.end

magic
tech gf180mcuD
magscale 1 10
timestamp 1755878577
<< polysilicon >>
rect 454 -742 514 -470
rect 618 -500 678 -470
rect 618 -560 839 -500
rect 779 -630 839 -560
rect 914 -574 1030 -514
rect 562 -698 678 -638
rect 779 -690 974 -630
rect 914 -741 974 -690
rect 1078 -742 1138 -470
rect 1374 -742 1434 -470
<< metal1 >>
rect 280 0 1772 140
rect 379 -143 425 0
rect 538 -698 562 -638
rect 622 -698 646 -638
rect 379 -980 425 -899
rect 707 -910 753 -132
rect 839 -910 885 -132
rect 1167 -143 1213 0
rect 1299 -143 1345 0
rect 946 -574 970 -514
rect 1030 -574 1054 -514
rect 1627 -630 1673 -457
rect 1463 -676 1673 -630
rect 1463 -755 1509 -676
rect 1167 -980 1213 -899
rect 1299 -980 1345 -899
rect 1627 -980 1673 -899
rect 280 -1120 1772 -980
<< via1 >>
rect 562 -698 622 -638
rect 970 -574 1030 -514
<< metal2 >>
rect 968 -514 1032 -496
rect 968 -570 970 -514
rect 560 -574 970 -570
rect 1030 -574 1032 -514
rect 560 -630 1032 -574
rect 560 -638 624 -630
rect 560 -698 562 -638
rect 622 -698 624 -638
rect 560 -716 624 -698
use nfet_03v3_C8ZVHP  nfet_03v3_C8ZVHP_0
timestamp 1755878577
transform 1 0 566 0 1 -827
box -224 -153 224 153
use nfet_03v3_C8ZVHP  nfet_03v3_C8ZVHP_1
timestamp 1755878577
transform 1 0 1026 0 1 -827
box -224 -153 224 153
use nfet_03v3_C8ZVHP  nfet_03v3_C8ZVHP_2
timestamp 1755878577
transform 1 0 1486 0 1 -827
box -224 -153 224 153
use pfet_03v3_XSR2S3  pfet_03v3_XSR2S3_0
timestamp 1755878577
transform -1 0 1486 0 1 -300
box -286 -300 286 300
use pfet_03v3_XSR2S3  pfet_03v3_XSR2S3_1
timestamp 1755878577
transform -1 0 1026 0 1 -300
box -286 -300 286 300
use pfet_03v3_XSR2S3  pfet_03v3_XSR2S3_2
timestamp 1755878577
transform -1 0 566 0 1 -300
box -286 -300 286 300
<< end >>

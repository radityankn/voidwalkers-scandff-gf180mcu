** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/schematics/mux2x1_transmission_gate/mux_toplevel.sch
.subckt mux_toplevel vdd data vss out scan_data se_in
*.PININFO vdd:B out:O data:I scan_data:I se_in:I vdd:B vss:B vss:B vdd:B vss:B
x2 vdd net1 data out se_in vss mux_tg
x3 vdd se_in scan_data out net1 vss mux_tg
x1 vdd se_in net1 vss mux_ctrl_logic
.ends

* expanding   symbol:  schematics/mux2x1_transmission_gate/mux_tg.sym # of pins=6
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/schematics/mux2x1_transmission_gate/mux_tg.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/schematics/mux2x1_transmission_gate/mux_tg.sch
.subckt mux_tg vdd pfet_gate in out nfet_gate gnd
*.PININFO vdd:B gnd:B out:B in:B pfet_gate:B nfet_gate:B
M1 in nfet_gate out gnd nfet_03v3 L=0.28u W=0.22u nf=1 m=1
M2 in pfet_gate out vdd pfet_03v3 L=0.28u W=0.22u nf=1 m=1
.ends


* expanding   symbol:  schematics/mux2x1_transmission_gate/mux_ctrl_logic.sym # of pins=4
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/schematics/mux2x1_transmission_gate/mux_ctrl_logic.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/schematics/mux2x1_transmission_gate/mux_ctrl_logic.sch
.subckt mux_ctrl_logic vdd in out_inv gnd
*.PININFO vdd:B gnd:B out_inv:B in:B
M1 out_inv in gnd gnd nfet_03v3 L=0.28u W=0.22u nf=1 m=1
M2 out_inv in vdd vdd pfet_03v3 L=0.28u W=0.22u nf=1 m=1
.ends


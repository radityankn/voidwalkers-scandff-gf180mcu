magic
tech gf180mcuD
magscale 1 10
timestamp 1756235029
<< nwell >>
rect 662 619 710 630
rect 1296 261 1302 265
rect 1296 249 1309 261
rect 1302 246 1309 249
rect 1311 246 1383 261
rect 1292 188 1643 246
rect 1302 182 1309 188
rect 1311 181 1383 188
<< pdiff >>
rect 662 619 710 630
<< ndiffc >>
rect 663 -195 709 -51
rect 991 -195 1037 -51
rect 1155 -195 1201 -51
rect 1319 -195 1365 -51
<< pdiffc >>
rect 663 305 709 619
rect 991 305 1037 619
rect 1319 305 1365 619
<< polysilicon >>
rect 323 735 634 795
rect 574 676 634 735
rect 410 266 470 315
rect 410 247 510 266
rect 410 187 430 247
rect 490 187 510 247
rect 410 166 510 187
rect 410 -45 470 166
rect 738 113 798 269
rect 862 248 962 270
rect 862 188 884 248
rect 944 188 962 248
rect 862 170 962 188
rect 518 69 798 113
rect 518 9 532 69
rect 592 54 798 69
rect 592 9 634 54
rect 518 -14 634 9
rect 902 6 962 170
rect 1066 161 1126 255
rect 1013 139 1126 161
rect 1013 79 1036 139
rect 1096 79 1126 139
rect 1013 59 1126 79
rect 1066 0 1126 59
rect 1230 134 1290 255
rect 1522 230 1637 257
rect 1522 179 1572 230
rect 1624 179 1637 230
rect 1522 158 1637 179
rect 1230 114 1350 134
rect 1230 54 1269 114
rect 1329 54 1350 114
rect 1230 34 1350 54
rect 1230 -41 1290 34
rect 1522 -2 1582 158
rect 1686 86 1746 262
rect 1632 65 1746 86
rect 1632 14 1651 65
rect 1703 14 1746 65
rect 1632 -6 1746 14
rect 1632 -7 1686 -6
rect 738 -312 798 -252
rect 333 -372 798 -312
<< polycontact >>
rect 430 187 490 247
rect 884 188 944 248
rect 532 9 592 69
rect 1036 79 1096 139
rect 1572 179 1624 230
rect 1269 54 1329 114
rect 1651 14 1703 65
<< metal1 >>
rect 236 706 1926 847
rect 334 303 382 706
rect 662 619 710 630
rect 662 305 663 619
rect 709 305 710 619
rect 410 187 430 247
rect 490 187 510 247
rect 662 139 710 305
rect 990 619 1038 706
rect 990 305 991 619
rect 1037 305 1038 619
rect 990 294 1038 305
rect 1318 619 1366 630
rect 1318 305 1319 619
rect 1365 305 1366 619
rect 1318 261 1366 305
rect 1302 248 1383 261
rect 862 188 884 248
rect 944 188 1314 248
rect 1374 246 1383 248
rect 1447 246 1493 302
rect 1611 294 1658 706
rect 1374 230 1643 246
rect 1374 188 1572 230
rect 662 138 751 139
rect 662 80 677 138
rect 735 80 751 138
rect 662 79 751 80
rect 1007 79 1036 139
rect 1096 79 1107 139
rect 513 9 532 69
rect 592 9 615 69
rect 334 -282 382 -41
rect 662 -51 710 79
rect 662 -195 663 -51
rect 709 -195 710 -51
rect 662 -206 710 -195
rect 990 -51 1038 -40
rect 990 -195 991 -51
rect 1037 -195 1038 -51
rect 990 -282 1038 -195
rect 1155 -51 1201 188
rect 1302 181 1383 188
rect 1248 54 1269 114
rect 1329 54 1348 114
rect 1447 70 1493 188
rect 1545 179 1572 188
rect 1624 179 1643 230
rect 1545 175 1643 179
rect 1775 165 1821 313
rect 1447 65 1725 70
rect 1447 14 1651 65
rect 1703 14 1725 65
rect 1447 10 1725 14
rect 1775 69 1932 165
rect 1155 -206 1201 -195
rect 1318 -51 1366 -28
rect 1447 -45 1493 10
rect 1318 -195 1319 -51
rect 1365 -195 1366 -51
rect 1318 -282 1366 -195
rect 1610 -282 1657 -41
rect 1775 -206 1821 69
rect 236 -423 1926 -282
<< via1 >>
rect 1314 188 1374 248
rect 677 80 735 138
<< metal2 >>
rect 1085 411 1223 471
rect 410 178 510 258
rect 677 142 735 150
rect 675 139 737 142
rect 1024 139 1107 149
rect 671 138 1107 139
rect 671 80 677 138
rect 735 80 1107 138
rect 513 0 614 80
rect 671 79 1107 80
rect 675 77 737 79
rect 677 68 735 77
rect 1024 69 1107 79
rect 1163 124 1223 411
rect 1302 248 1383 261
rect 1302 188 1314 248
rect 1374 246 1383 248
rect 1374 243 1643 246
rect 1374 188 1646 243
rect 1302 182 1383 188
rect 1303 181 1383 182
rect 1546 168 1646 188
rect 1163 54 1349 124
rect 1179 53 1349 54
rect 1237 45 1349 53
rect 533 -81 593 0
rect 236 -141 593 -81
use nfet_03v3_C8ZVHP  nfet_03v3_C8ZVHP_0
timestamp 1756212155
transform 1 0 1634 0 1 -123
box -200 -129 200 129
use nfet_03v3_CYXVHP  nfet_03v3_CYXVHP_0
timestamp 1756235029
transform 1 0 850 0 1 -123
box -528 -129 528 129
use pfet_03v3_XSR2S3  pfet_03v3_XSR2S3_0
timestamp 1756212155
transform 1 0 1634 0 1 462
box -286 -300 286 300
use pfet_03v3_XSV2S3  pfet_03v3_XSV2S3_0
timestamp 1756235029
transform 1 0 850 0 1 462
box -614 -300 614 300
<< end >>

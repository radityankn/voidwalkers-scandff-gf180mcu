magic
tech gf180mcuD
magscale 1 10
timestamp 1756653248
<< error_s >>
rect -960 340 -957 470
<< nwell >>
rect -970 650 2610 1370
<< pwell >>
rect -970 540 2610 650
rect -970 520 1960 540
rect 2090 520 2150 540
rect 2280 520 2340 540
rect 2420 520 2610 540
rect -970 100 2610 520
<< nmos >>
rect -870 320 -810 490
rect -680 320 -620 490
rect -490 320 -430 490
rect -340 320 -280 490
rect 10 320 70 490
rect 120 320 180 490
rect 310 320 370 490
rect 790 320 850 490
rect 1180 320 1240 490
rect 1370 320 1430 490
rect 1560 320 1620 490
rect 1710 320 1770 490
rect 1900 320 1960 490
rect 2090 320 2150 490
rect 2280 320 2340 490
<< pmos >>
rect -840 810 -780 1150
rect -730 810 -670 1150
rect -490 810 -430 1150
rect -340 810 -280 1150
rect -150 810 -90 1150
rect 120 810 180 1150
rect 310 810 370 1150
rect 790 810 850 1150
rect 1210 810 1270 1150
rect 1370 810 1430 1150
rect 1560 810 1620 1150
rect 1710 810 1770 1150
rect 1900 810 1960 1150
rect 2090 810 2150 1150
rect 2280 810 2340 1150
<< ndiff >>
rect -970 470 -870 490
rect -970 340 -960 470
rect -910 340 -870 470
rect -970 320 -870 340
rect -810 470 -680 490
rect -810 340 -780 470
rect -710 340 -680 470
rect -810 320 -680 340
rect -620 450 -490 490
rect -620 340 -580 450
rect -530 340 -490 450
rect -620 320 -490 340
rect -430 320 -340 490
rect -280 430 10 490
rect -280 340 -250 430
rect -200 340 10 430
rect -280 320 10 340
rect 70 320 120 490
rect 180 400 310 490
rect 180 340 220 400
rect 270 340 310 400
rect 180 320 310 340
rect 370 470 550 490
rect 370 340 410 470
rect 460 340 550 470
rect 370 320 550 340
rect 680 470 790 490
rect 680 340 700 470
rect 750 340 790 470
rect 680 320 790 340
rect 850 470 1000 490
rect 850 340 930 470
rect 980 340 1000 470
rect 850 320 1000 340
rect 1070 470 1180 490
rect 1070 340 1090 470
rect 1140 340 1180 470
rect 1070 320 1180 340
rect 1240 470 1370 490
rect 1240 340 1270 470
rect 1340 340 1370 470
rect 1240 320 1370 340
rect 1430 470 1560 490
rect 1430 340 1470 470
rect 1520 340 1560 470
rect 1430 320 1560 340
rect 1620 320 1710 490
rect 1770 470 1900 490
rect 1770 340 1810 470
rect 1860 340 1900 470
rect 1770 320 1900 340
rect 1960 320 2090 490
rect 2150 470 2280 490
rect 2150 340 2190 470
rect 2240 340 2280 470
rect 2150 320 2280 340
rect 2340 470 2520 490
rect 2340 340 2380 470
rect 2430 340 2520 470
rect 2340 320 2520 340
<< pdiff >>
rect -950 1130 -840 1150
rect -950 1010 -930 1130
rect -880 1010 -840 1130
rect -950 950 -840 1010
rect -950 830 -930 950
rect -880 830 -840 950
rect -950 810 -840 830
rect -780 810 -730 1150
rect -670 1130 -490 1150
rect -670 1010 -610 1130
rect -560 1010 -490 1130
rect -670 810 -490 1010
rect -430 810 -340 1150
rect -280 1130 -150 1150
rect -280 1010 -250 1130
rect -200 1010 -150 1130
rect -280 810 -150 1010
rect -90 810 120 1150
rect 180 1130 310 1150
rect 180 1010 220 1130
rect 270 1010 310 1130
rect 180 810 310 1010
rect 370 950 550 1150
rect 370 830 460 950
rect 510 830 550 950
rect 370 810 550 830
rect 680 1130 790 1150
rect 680 1010 700 1130
rect 750 1010 790 1130
rect 680 810 790 1010
rect 850 950 1000 1150
rect 850 830 930 950
rect 980 830 1000 950
rect 850 810 1000 830
rect 1100 1130 1210 1150
rect 1100 1010 1120 1130
rect 1170 1010 1210 1130
rect 1100 950 1210 1010
rect 1100 830 1120 950
rect 1170 830 1210 950
rect 1100 810 1210 830
rect 1270 810 1370 1150
rect 1430 1130 1560 1150
rect 1430 1010 1470 1130
rect 1520 1010 1560 1130
rect 1430 950 1560 1010
rect 1430 830 1470 950
rect 1520 830 1560 950
rect 1430 810 1560 830
rect 1620 810 1710 1150
rect 1770 1130 1900 1150
rect 1770 1010 1810 1130
rect 1860 1010 1900 1130
rect 1770 950 1900 1010
rect 1770 830 1810 950
rect 1860 830 1900 950
rect 1770 810 1900 830
rect 1960 810 2090 1150
rect 2150 1130 2280 1150
rect 2150 1010 2190 1130
rect 2240 1010 2280 1130
rect 2150 950 2280 1010
rect 2150 830 2190 950
rect 2240 830 2280 950
rect 2150 810 2280 830
rect 2340 950 2520 1150
rect 2340 830 2430 950
rect 2480 830 2520 950
rect 2340 810 2520 830
<< ndiffc >>
rect -960 340 -910 470
rect -780 340 -710 470
rect -580 340 -530 450
rect -250 340 -200 430
rect 220 340 270 400
rect 410 340 460 470
rect 700 340 750 470
rect 930 340 980 470
rect 1090 340 1140 470
rect 1270 340 1340 470
rect 1470 340 1520 470
rect 1810 340 1860 470
rect 2190 340 2240 470
rect 2380 340 2430 470
<< pdiffc >>
rect -930 1010 -880 1130
rect -930 830 -880 950
rect -610 1010 -560 1130
rect -250 1010 -200 1130
rect 220 1010 270 1130
rect 460 830 510 950
rect 700 1010 750 1130
rect 930 830 980 950
rect 1120 1010 1170 1130
rect 1120 830 1170 950
rect 1470 1010 1520 1130
rect 1470 830 1520 950
rect 1810 1010 1860 1130
rect 1810 830 1860 950
rect 2190 1010 2240 1130
rect 2190 830 2240 950
rect 2430 830 2480 950
<< polysilicon >>
rect -840 1250 850 1310
rect -840 1150 -780 1250
rect -730 1150 -670 1200
rect -490 1150 -430 1200
rect -340 1150 -280 1200
rect -150 1150 -90 1200
rect 120 1150 180 1200
rect 310 1150 370 1200
rect 790 1150 850 1250
rect 1900 1250 2340 1310
rect 1210 1150 1270 1200
rect 1370 1150 1430 1200
rect 1560 1150 1620 1200
rect 1710 1150 1770 1200
rect 1900 1150 1960 1250
rect 2090 1150 2150 1200
rect 2280 1150 2340 1250
rect -840 780 -780 810
rect -870 660 -780 780
rect -730 780 -670 810
rect -490 780 -430 810
rect -730 760 -620 780
rect -730 690 -710 760
rect -640 690 -620 760
rect -730 670 -620 690
rect -560 720 -430 780
rect -340 780 -280 810
rect -340 760 -240 780
rect -150 760 -90 810
rect 120 780 180 810
rect 120 760 240 780
rect -870 490 -810 660
rect -730 580 -670 670
rect -560 610 -490 720
rect -340 680 -320 760
rect -260 680 -240 760
rect -340 660 -240 680
rect -170 740 -70 760
rect -170 650 -150 740
rect -90 650 -70 740
rect -170 630 -70 650
rect -20 740 70 760
rect -20 670 0 740
rect 50 670 70 740
rect -560 590 -430 610
rect -730 520 -620 580
rect -560 540 -540 590
rect -490 540 -430 590
rect -150 580 -90 630
rect -560 520 -430 540
rect -680 490 -620 520
rect -490 490 -430 520
rect -340 520 -90 580
rect -20 540 70 670
rect -340 490 -280 520
rect 10 490 70 540
rect 120 700 140 760
rect 220 700 240 760
rect 120 680 240 700
rect 120 490 180 680
rect 310 490 370 810
rect 790 490 850 810
rect 1210 780 1270 810
rect 1110 760 1270 780
rect 1110 680 1130 760
rect 1220 680 1270 760
rect 1110 660 1270 680
rect 1370 780 1430 810
rect 1370 760 1510 780
rect 1370 690 1420 760
rect 1490 690 1510 760
rect 1370 670 1510 690
rect 1180 490 1240 660
rect 1370 490 1430 670
rect 1560 650 1620 810
rect 1710 710 1770 810
rect 1900 760 1960 810
rect 2090 780 2150 810
rect 2090 760 2210 780
rect 1710 650 1960 710
rect 1560 630 1660 650
rect 1560 560 1580 630
rect 1640 560 1660 630
rect 1560 540 1660 560
rect 1900 630 1960 650
rect 2090 700 2110 760
rect 2190 700 2210 760
rect 2090 680 2210 700
rect 2280 700 2340 810
rect 1900 610 2020 630
rect 1900 560 1920 610
rect 2000 560 2020 610
rect 1900 540 2020 560
rect 1560 490 1620 540
rect 1710 490 1770 540
rect 1900 490 1960 540
rect 2090 490 2150 680
rect 2280 640 2580 700
rect 2280 490 2340 640
rect -870 270 -810 320
rect -680 270 -620 320
rect -490 270 -430 320
rect -340 270 -280 320
rect 10 220 70 320
rect 120 270 180 320
rect 310 220 370 320
rect 790 270 850 320
rect 1180 270 1240 320
rect 1370 270 1430 320
rect 1560 270 1620 320
rect 1710 220 1770 320
rect 1900 270 1960 320
rect 2090 270 2150 320
rect 2280 220 2340 320
rect 10 160 2340 220
<< polycontact >>
rect -710 690 -640 760
rect -320 680 -260 760
rect -150 650 -90 740
rect 0 670 50 740
rect -540 540 -490 590
rect 140 700 220 760
rect 1130 680 1220 760
rect 1420 690 1490 760
rect 1580 560 1640 630
rect 2110 700 2190 760
rect 1920 560 2000 610
<< metal1 >>
rect -970 1250 2610 1370
rect -970 1130 -870 1150
rect -970 1020 -930 1130
rect -940 1010 -930 1020
rect -880 1010 -870 1130
rect -940 950 -870 1010
rect -620 1130 -550 1250
rect -620 1010 -610 1130
rect -560 1010 -550 1130
rect -620 990 -550 1010
rect -500 1130 -180 1150
rect -500 1010 -250 1130
rect -200 1010 -180 1130
rect -500 990 -180 1010
rect 210 1130 280 1250
rect 210 1010 220 1130
rect 270 1010 280 1130
rect 210 990 280 1010
rect 330 1020 640 1150
rect -940 830 -930 950
rect -880 830 -870 950
rect -500 940 -440 990
rect 330 940 400 1020
rect -940 610 -870 830
rect -730 880 -440 940
rect -730 760 -620 880
rect -730 690 -710 760
rect -640 720 -620 760
rect -340 820 70 940
rect -340 760 -240 820
rect -640 690 -390 720
rect -730 660 -390 690
rect -340 680 -320 760
rect -260 680 -240 760
rect -340 660 -240 680
rect -150 740 -70 760
rect -940 590 -490 610
rect -940 540 -540 590
rect -780 520 -490 540
rect -970 470 -900 490
rect -970 340 -960 470
rect -910 340 -900 470
rect -970 220 -900 340
rect -780 470 -700 520
rect -710 340 -700 470
rect -780 320 -700 340
rect -590 450 -520 470
rect -590 340 -580 450
rect -530 340 -520 450
rect -590 220 -520 340
rect -440 430 -390 660
rect -90 650 -70 740
rect -150 530 -70 650
rect 0 740 70 820
rect 50 670 70 740
rect 120 880 400 940
rect 450 950 520 970
rect 120 760 240 880
rect 120 700 140 760
rect 220 700 240 760
rect 450 830 460 950
rect 510 830 520 950
rect 570 940 640 1020
rect 690 1130 760 1250
rect 690 1010 700 1130
rect 750 1010 760 1130
rect 690 990 760 1010
rect 810 1130 1350 1150
rect 810 1020 1120 1130
rect 810 940 870 1020
rect 1110 1010 1120 1020
rect 1170 1030 1350 1130
rect 1170 1010 1180 1030
rect 570 870 870 940
rect 920 950 1060 970
rect 0 580 70 670
rect 450 530 520 830
rect 920 830 930 950
rect 980 830 1060 950
rect 920 810 1060 830
rect 1110 950 1180 1010
rect 1110 830 1120 950
rect 1170 830 1180 950
rect 1110 810 1180 830
rect 1000 760 1060 810
rect 1000 680 1130 760
rect 1220 680 1240 760
rect 1000 610 1060 680
rect -150 470 520 530
rect 920 540 1060 610
rect 1290 630 1350 1030
rect 1460 1130 1530 1250
rect 1460 1010 1470 1130
rect 1520 1010 1530 1130
rect 1460 950 1530 1010
rect 1460 830 1470 950
rect 1520 830 1530 950
rect 1460 810 1530 830
rect 1580 1130 1870 1150
rect 1580 1030 1810 1130
rect 1580 760 1650 1030
rect 1400 690 1420 760
rect 1490 690 1650 760
rect 1400 680 1650 690
rect 1800 1010 1810 1030
rect 1860 1010 1870 1130
rect 1800 950 1870 1010
rect 1800 830 1810 950
rect 1860 830 1870 950
rect 1290 560 1580 630
rect 1640 560 1660 630
rect 1290 540 1660 560
rect -440 340 -250 430
rect -200 340 -180 430
rect -440 320 -180 340
rect 210 400 280 420
rect 210 340 220 400
rect 270 340 280 400
rect 210 220 280 340
rect 400 340 410 470
rect 460 340 520 470
rect 400 320 520 340
rect 690 470 760 490
rect 690 340 700 470
rect 750 340 760 470
rect 690 220 760 340
rect 920 470 990 540
rect 1290 490 1350 540
rect 920 340 930 470
rect 980 340 990 470
rect 920 320 990 340
rect 1080 470 1150 490
rect 1080 340 1090 470
rect 1140 340 1150 470
rect 1080 220 1150 340
rect 1270 470 1350 490
rect 1340 340 1350 470
rect 1270 320 1350 340
rect 1460 470 1530 490
rect 1460 340 1470 470
rect 1520 340 1530 470
rect 1460 220 1530 340
rect 1800 470 1870 830
rect 2180 1130 2250 1250
rect 2180 1010 2190 1130
rect 2240 1010 2250 1130
rect 2180 950 2250 1010
rect 2180 830 2190 950
rect 2240 830 2250 950
rect 2180 810 2250 830
rect 2300 1020 2610 1150
rect 2300 760 2370 1020
rect 2090 700 2110 760
rect 2190 700 2370 760
rect 2420 950 2490 970
rect 2420 830 2430 950
rect 2480 830 2490 950
rect 2420 630 2490 830
rect 1920 610 2490 630
rect 2000 560 2490 610
rect 1920 540 2490 560
rect 2420 490 2490 540
rect 1800 340 1810 470
rect 1860 340 1870 470
rect 1800 320 1870 340
rect 2180 470 2250 490
rect 2180 340 2190 470
rect 2240 340 2250 470
rect 2180 220 2250 340
rect 2370 470 2490 490
rect 2370 340 2380 470
rect 2430 340 2490 470
rect 2370 320 2490 340
rect -970 100 2610 220
use inverter_component  inverter_component_0
timestamp 1756652194
transform 1 0 -1420 0 1 350
box -260 -250 450 1020
use mux_component  mux_component_0
timestamp 1756653248
transform 1 0 2280 0 1 350
box 330 -250 1510 1020
<< end >>

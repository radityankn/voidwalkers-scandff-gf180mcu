magic
tech gf180mcuD
magscale 1 10
timestamp 1755874087
<< nwell >>
rect 96 138 144 468
rect 260 132 308 548
rect 916 132 964 556
rect 172 1 282 88
rect 172 0 232 1
rect 1274 0 2666 600
<< pwell >>
rect -6 -462 2670 0
<< nmos >>
rect 1448 -380 1508 -210
rect 1612 -380 1672 -210
rect 1776 -380 1836 -210
rect 1940 -380 2000 -210
rect 2104 -380 2164 -210
rect 2268 -380 2328 -210
rect 2432 -380 2492 -210
<< pmos >>
rect 1448 130 1508 470
rect 1612 130 1672 470
rect 1776 130 1836 470
rect 1940 130 2000 470
rect 2104 130 2164 470
rect 2268 130 2328 470
rect 2432 130 2492 470
<< ndiff >>
rect 1360 -223 1448 -210
rect 1360 -367 1373 -223
rect 1419 -367 1448 -223
rect 1360 -380 1448 -367
rect 1508 -223 1612 -210
rect 1508 -367 1537 -223
rect 1583 -367 1612 -223
rect 1508 -380 1612 -367
rect 1672 -223 1776 -210
rect 1672 -367 1701 -223
rect 1747 -367 1776 -223
rect 1672 -380 1776 -367
rect 1836 -223 1940 -210
rect 1836 -367 1865 -223
rect 1911 -367 1940 -223
rect 1836 -380 1940 -367
rect 2000 -223 2104 -210
rect 2000 -367 2029 -223
rect 2075 -367 2104 -223
rect 2000 -380 2104 -367
rect 2164 -223 2268 -210
rect 2164 -367 2193 -223
rect 2239 -367 2268 -223
rect 2164 -380 2268 -367
rect 2328 -223 2432 -210
rect 2328 -367 2357 -223
rect 2403 -367 2432 -223
rect 2328 -380 2432 -367
rect 2492 -223 2580 -210
rect 2492 -367 2521 -223
rect 2567 -367 2580 -223
rect 2492 -380 2580 -367
<< pdiff >>
rect 1360 457 1448 470
rect 1360 143 1373 457
rect 1419 143 1448 457
rect 1360 130 1448 143
rect 1508 457 1612 470
rect 1508 143 1537 457
rect 1583 143 1612 457
rect 1508 130 1612 143
rect 1672 457 1776 470
rect 1672 143 1701 457
rect 1747 143 1776 457
rect 1672 130 1776 143
rect 1836 457 1940 470
rect 1836 143 1865 457
rect 1911 143 1940 457
rect 1836 130 1940 143
rect 2000 457 2104 470
rect 2000 143 2029 457
rect 2075 143 2104 457
rect 2000 130 2104 143
rect 2164 457 2268 470
rect 2164 143 2193 457
rect 2239 143 2268 457
rect 2164 130 2268 143
rect 2328 457 2432 470
rect 2328 143 2357 457
rect 2403 143 2432 457
rect 2328 130 2432 143
rect 2492 457 2580 470
rect 2492 143 2521 457
rect 2567 143 2580 457
rect 2492 130 2580 143
<< ndiffc >>
rect 1373 -367 1419 -223
rect 1537 -367 1583 -223
rect 1701 -367 1747 -223
rect 1865 -367 1911 -223
rect 2029 -367 2075 -223
rect 2193 -367 2239 -223
rect 2357 -367 2403 -223
rect 2521 -367 2567 -223
<< pdiffc >>
rect 1373 143 1419 457
rect 1537 143 1583 457
rect 1701 143 1747 457
rect 1865 143 1911 457
rect 2029 143 2075 457
rect 2193 143 2239 457
rect 2357 143 2403 457
rect 2521 143 2567 457
<< polysilicon >>
rect 1448 470 1508 514
rect 1612 470 1672 514
rect 1776 470 1836 514
rect 1940 470 2000 514
rect 2104 470 2164 514
rect 2268 470 2328 514
rect 2432 470 2492 514
rect 172 74 282 88
rect 172 14 207 74
rect 267 14 282 74
rect 172 1 282 14
rect 172 -206 232 1
rect 336 -166 396 86
rect 828 -166 888 86
rect 992 0 1052 86
rect 969 -21 1069 0
rect 969 -81 990 -21
rect 1050 -81 1069 -21
rect 969 -100 1069 -81
rect 992 -166 1052 -100
rect 1156 -170 1216 86
rect 1448 -210 1508 130
rect 1612 0 1672 130
rect 1595 -21 1695 0
rect 1595 -81 1614 -21
rect 1674 -81 1695 -21
rect 1595 -100 1695 -81
rect 1612 -210 1672 -100
rect 1776 -210 1836 130
rect 1940 86 2000 130
rect 2104 86 2164 130
rect 1940 -210 2000 -166
rect 2104 -210 2164 -166
rect 2268 -210 2328 130
rect 2432 88 2492 130
rect 2382 74 2492 88
rect 2382 14 2397 74
rect 2457 14 2492 74
rect 2382 1 2492 14
rect 2432 -210 2492 1
rect 1448 -424 1508 -380
rect 1612 -424 1672 -380
rect 1776 -424 1836 -380
rect 1940 -424 2000 -380
rect 2104 -424 2164 -380
rect 2268 -424 2328 -380
rect 2432 -424 2492 -380
<< polycontact >>
rect 207 14 267 74
rect 990 -81 1050 -21
rect 1614 -81 1674 -21
rect 2397 14 2457 74
<< metal1 >>
rect -2 544 2666 684
rect 96 -110 144 468
rect 260 132 308 544
rect 196 74 278 85
rect 196 14 207 74
rect 267 14 278 74
rect 196 3 278 14
rect 588 -7 636 468
rect 916 132 964 544
rect 1373 457 1419 468
rect 1373 132 1419 143
rect 1537 457 1583 468
rect 1537 132 1583 143
rect 1700 457 1748 544
rect 1700 143 1701 457
rect 1747 143 1748 457
rect 1700 132 1748 143
rect 1865 457 1911 468
rect 1865 132 1911 143
rect 2028 457 2076 468
rect 2028 143 2029 457
rect 2075 143 2076 457
rect 2028 -7 2076 143
rect 2193 457 2239 468
rect 2193 132 2239 143
rect 2356 457 2404 544
rect 2356 143 2357 457
rect 2403 143 2404 457
rect 2356 132 2404 143
rect 2520 457 2568 468
rect 2520 143 2521 457
rect 2567 143 2568 457
rect 2386 74 2468 85
rect 2386 14 2397 74
rect 2457 14 2468 74
rect 2386 3 2468 14
rect 570 -18 654 -7
rect 570 -78 582 -18
rect 642 -20 654 -18
rect 977 -20 1062 -8
rect 642 -21 1062 -20
rect 642 -78 990 -21
rect 570 -91 654 -78
rect 977 -81 990 -78
rect 1050 -81 1062 -21
rect 78 -122 162 -110
rect 78 -182 90 -122
rect 150 -182 162 -122
rect 78 -194 162 -182
rect 96 -372 144 -194
rect 260 -454 308 -204
rect 588 -370 636 -91
rect 977 -93 1062 -81
rect 1602 -20 1687 -8
rect 2010 -18 2094 -7
rect 2010 -20 2022 -18
rect 1602 -21 2022 -20
rect 1602 -81 1614 -21
rect 1674 -78 2022 -21
rect 2082 -78 2094 -18
rect 1674 -81 1687 -78
rect 1602 -93 1687 -81
rect 2010 -91 2094 -78
rect 916 -454 964 -204
rect 1244 -454 1292 -204
rect 1372 -223 1420 -204
rect 1372 -367 1373 -223
rect 1419 -367 1420 -223
rect 1372 -454 1420 -367
rect 1537 -223 1583 -212
rect 1537 -378 1583 -367
rect 1700 -223 1748 -204
rect 1700 -367 1701 -223
rect 1747 -367 1748 -223
rect 1700 -454 1748 -367
rect 1865 -223 1911 -212
rect 1865 -378 1911 -367
rect 2028 -223 2076 -91
rect 2520 -110 2568 143
rect 2502 -122 2586 -110
rect 2502 -182 2514 -122
rect 2574 -182 2586 -122
rect 2502 -194 2586 -182
rect 2028 -367 2029 -223
rect 2075 -367 2076 -223
rect 2028 -370 2076 -367
rect 2193 -223 2239 -212
rect 2029 -378 2075 -370
rect 2193 -378 2239 -367
rect 2356 -223 2404 -204
rect 2356 -367 2357 -223
rect 2403 -367 2404 -223
rect 2356 -454 2404 -367
rect 2520 -223 2568 -194
rect 2520 -367 2521 -223
rect 2567 -367 2568 -223
rect 2520 -372 2568 -367
rect 2521 -378 2567 -372
rect -8 -594 2672 -454
<< via1 >>
rect 582 -78 642 -18
rect 90 -182 150 -122
rect 2022 -78 2082 -18
rect 2514 -182 2574 -122
<< metal2 >>
rect 570 -18 654 -7
rect 570 -78 582 -18
rect 642 -78 654 -18
rect 570 -91 654 -78
rect 2010 -18 2094 -7
rect 2010 -78 2022 -18
rect 2082 -78 2094 -18
rect 2010 -91 2094 -78
rect 78 -122 162 -110
rect 78 -182 90 -122
rect 150 -182 162 -122
rect 78 -194 162 -182
rect 2502 -122 2586 -110
rect 2502 -182 2514 -122
rect 2574 -182 2586 -122
rect 2502 -194 2586 -182
use nfet_03v3_CWXVHP  nfet_03v3_CWXVHP_0
timestamp 1755874087
transform 1 0 694 0 1 -295
box -610 -129 610 129
use nfet_03v3_CWXVHP  nfet_03v3_CWXVHP_1
timestamp 1755874087
transform -1 0 1970 0 1 -295
box -610 -129 610 129
use pfet_03v3_XSU2S3  pfet_03v3_XSU2S3_0
timestamp 1755830194
transform 1 0 694 0 1 300
box -696 -300 696 300
use pfet_03v3_XSU2S3  pfet_03v3_XSU2S3_1
timestamp 1755830194
transform -1 0 1970 0 1 300
box -696 -300 696 300
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1756740167
<< nwell >>
rect -1690 650 2660 1370
<< pwell >>
rect -1690 540 2660 650
rect -1690 520 1960 540
rect 2090 520 2150 540
rect 2280 520 2340 540
rect 2420 520 2660 540
rect -1690 100 2660 520
<< nmos >>
rect -1490 320 -1430 490
rect -1300 320 -1240 490
rect -870 320 -810 490
rect -680 320 -620 490
rect -490 320 -430 490
rect -340 320 -280 490
rect 10 320 70 490
rect 120 320 180 490
rect 310 320 370 490
rect 790 320 850 490
rect 1180 320 1240 490
rect 1370 320 1430 490
rect 1560 320 1620 490
rect 1710 320 1770 490
rect 1900 320 1960 490
rect 2090 320 2150 490
rect 2280 320 2340 490
<< pmos >>
rect -1490 810 -1430 1150
rect -1300 810 -1240 1150
rect -840 810 -780 1150
rect -730 810 -670 1150
rect -490 810 -430 1150
rect -340 810 -280 1150
rect -150 810 -90 1150
rect 120 810 180 1150
rect 310 810 370 1150
rect 790 800 850 1140
rect 1210 810 1270 1150
rect 1370 810 1430 1150
rect 1560 810 1620 1150
rect 1710 810 1770 1150
rect 1900 810 1960 1150
rect 2090 810 2150 1150
rect 2280 810 2340 1150
<< ndiff >>
rect -1600 428 -1490 490
rect -1600 382 -1578 428
rect -1532 382 -1490 428
rect -1600 320 -1490 382
rect -1430 428 -1300 490
rect -1430 382 -1388 428
rect -1342 382 -1300 428
rect -1430 320 -1300 382
rect -1240 428 -1111 490
rect -1240 382 -1198 428
rect -1152 382 -1111 428
rect -1240 320 -1111 382
rect -980 428 -870 490
rect -980 382 -958 428
rect -912 382 -870 428
rect -980 320 -870 382
rect -810 428 -680 490
rect -810 382 -768 428
rect -722 382 -680 428
rect -810 320 -680 382
rect -620 418 -490 490
rect -620 372 -578 418
rect -532 372 -490 418
rect -620 320 -490 372
rect -430 320 -340 490
rect -280 408 10 490
rect -280 362 -248 408
rect -202 362 10 408
rect -280 320 10 362
rect 70 320 120 490
rect 180 393 310 490
rect 180 347 222 393
rect 268 347 310 393
rect 180 320 310 347
rect 370 428 550 490
rect 370 382 412 428
rect 458 382 550 428
rect 370 320 550 382
rect 680 428 790 490
rect 680 382 702 428
rect 748 382 790 428
rect 680 320 790 382
rect 850 428 1000 490
rect 850 382 932 428
rect 978 382 1000 428
rect 850 320 1000 382
rect 1070 428 1180 490
rect 1070 382 1092 428
rect 1138 382 1180 428
rect 1070 320 1180 382
rect 1240 428 1370 490
rect 1240 382 1282 428
rect 1328 382 1370 428
rect 1240 320 1370 382
rect 1430 428 1560 490
rect 1430 382 1472 428
rect 1518 382 1560 428
rect 1430 320 1560 382
rect 1620 320 1710 490
rect 1770 428 1900 490
rect 1770 382 1812 428
rect 1858 382 1900 428
rect 1770 320 1900 382
rect 1960 320 2090 490
rect 2150 428 2280 490
rect 2150 382 2192 428
rect 2238 382 2280 428
rect 2150 320 2280 382
rect 2340 428 2520 490
rect 2340 382 2382 428
rect 2428 382 2520 428
rect 2340 320 2520 382
<< pdiff >>
rect -1600 1093 -1490 1150
rect -1600 1047 -1578 1093
rect -1532 1047 -1490 1093
rect -1600 810 -1490 1047
rect -1430 1093 -1300 1150
rect -1430 1047 -1388 1093
rect -1342 1047 -1300 1093
rect -1430 913 -1300 1047
rect -1430 867 -1388 913
rect -1342 867 -1300 913
rect -1430 810 -1300 867
rect -1240 1093 -1111 1150
rect -1240 1047 -1198 1093
rect -1152 1047 -1111 1093
rect -1240 913 -1111 1047
rect -1240 867 -1198 913
rect -1152 867 -1111 913
rect -1240 810 -1111 867
rect -950 1093 -840 1150
rect -950 1047 -928 1093
rect -882 1047 -840 1093
rect -950 913 -840 1047
rect -950 867 -928 913
rect -882 867 -840 913
rect -950 810 -840 867
rect -780 810 -730 1150
rect -670 1093 -490 1150
rect -670 1047 -608 1093
rect -562 1047 -490 1093
rect -670 810 -490 1047
rect -430 810 -340 1150
rect -280 1093 -150 1150
rect -280 1047 -248 1093
rect -202 1047 -150 1093
rect -280 810 -150 1047
rect -90 810 120 1150
rect 180 1093 310 1150
rect 180 1047 222 1093
rect 268 1047 310 1093
rect 180 810 310 1047
rect 370 913 550 1150
rect 370 867 462 913
rect 508 867 550 913
rect 370 810 550 867
rect 680 1083 790 1140
rect 680 1037 702 1083
rect 748 1037 790 1083
rect 680 800 790 1037
rect 850 913 1000 1140
rect 850 867 932 913
rect 978 867 1000 913
rect 850 800 1000 867
rect 1100 1093 1210 1150
rect 1100 1047 1122 1093
rect 1168 1047 1210 1093
rect 1100 913 1210 1047
rect 1100 867 1122 913
rect 1168 867 1210 913
rect 1100 810 1210 867
rect 1270 810 1370 1150
rect 1430 1093 1560 1150
rect 1430 1047 1472 1093
rect 1518 1047 1560 1093
rect 1430 913 1560 1047
rect 1430 867 1472 913
rect 1518 867 1560 913
rect 1430 810 1560 867
rect 1620 810 1710 1150
rect 1770 1093 1900 1150
rect 1770 1047 1812 1093
rect 1858 1047 1900 1093
rect 1770 913 1900 1047
rect 1770 867 1812 913
rect 1858 867 1900 913
rect 1770 810 1900 867
rect 1960 810 2090 1150
rect 2150 1093 2280 1150
rect 2150 1047 2192 1093
rect 2238 1047 2280 1093
rect 2150 913 2280 1047
rect 2150 867 2192 913
rect 2238 867 2280 913
rect 2150 810 2280 867
rect 2340 913 2520 1150
rect 2340 867 2432 913
rect 2478 867 2520 913
rect 2340 810 2520 867
<< ndiffc >>
rect -1578 382 -1532 428
rect -1388 382 -1342 428
rect -1198 382 -1152 428
rect -958 382 -912 428
rect -768 382 -722 428
rect -578 372 -532 418
rect -248 362 -202 408
rect 222 347 268 393
rect 412 382 458 428
rect 702 382 748 428
rect 932 382 978 428
rect 1092 382 1138 428
rect 1282 382 1328 428
rect 1472 382 1518 428
rect 1812 382 1858 428
rect 2192 382 2238 428
rect 2382 382 2428 428
<< pdiffc >>
rect -1578 1047 -1532 1093
rect -1388 1047 -1342 1093
rect -1388 867 -1342 913
rect -1198 1047 -1152 1093
rect -1198 867 -1152 913
rect -928 1047 -882 1093
rect -928 867 -882 913
rect -608 1047 -562 1093
rect -248 1047 -202 1093
rect 222 1047 268 1093
rect 462 867 508 913
rect 702 1037 748 1083
rect 932 867 978 913
rect 1122 1047 1168 1093
rect 1122 867 1168 913
rect 1472 1047 1518 1093
rect 1472 867 1518 913
rect 1812 1047 1858 1093
rect 1812 867 1858 913
rect 2192 1047 2238 1093
rect 2192 867 2238 913
rect 2432 867 2478 913
<< psubdiff >>
rect -1650 198 -1510 220
rect -1650 152 -1603 198
rect -1557 152 -1510 198
rect -1650 130 -1510 152
rect -880 198 -640 220
rect -880 152 -830 198
rect -690 152 -640 198
rect -880 130 -640 152
rect -270 198 -30 220
rect -270 152 -220 198
rect -80 152 -30 198
rect 2370 198 2610 220
rect -270 130 -30 152
rect 2370 152 2420 198
rect 2560 152 2610 198
rect 2370 130 2610 152
<< nsubdiff >>
rect -1600 1318 -1440 1340
rect -1600 1272 -1543 1318
rect -1497 1272 -1440 1318
rect -1600 1250 -1440 1272
rect 2370 1318 2610 1340
rect 600 1268 740 1290
rect 600 1222 647 1268
rect 693 1222 740 1268
rect 600 1200 740 1222
rect 2370 1272 2420 1318
rect 2560 1272 2610 1318
rect 2370 1250 2610 1272
<< psubdiffcont >>
rect -1603 152 -1557 198
rect -830 152 -690 198
rect -220 152 -80 198
rect 2420 152 2560 198
<< nsubdiffcont >>
rect -1543 1272 -1497 1318
rect 647 1222 693 1268
rect 2420 1272 2560 1318
<< polysilicon >>
rect -840 1310 1270 1350
rect -1490 1150 -1430 1200
rect -1300 1150 -1240 1200
rect -840 1150 -780 1310
rect -730 1150 -670 1200
rect -490 1150 -430 1200
rect -340 1150 -280 1200
rect -150 1150 -90 1200
rect 120 1150 180 1200
rect 310 1150 370 1200
rect 790 1140 850 1200
rect 1210 1150 1270 1310
rect 1900 1250 2340 1310
rect 1370 1150 1430 1200
rect 1560 1150 1620 1200
rect 1710 1150 1770 1200
rect 1900 1150 1960 1250
rect 2090 1150 2150 1200
rect 2280 1150 2340 1250
rect -1490 640 -1430 810
rect -1300 760 -1240 810
rect -840 780 -780 810
rect -1300 733 -990 760
rect -1300 687 -1073 733
rect -1027 687 -990 733
rect -1300 660 -990 687
rect -870 660 -780 780
rect -730 780 -670 810
rect -490 780 -430 810
rect -730 748 -620 780
rect -730 702 -698 748
rect -652 702 -620 748
rect -730 670 -620 702
rect -560 720 -430 780
rect -340 780 -280 810
rect -340 743 -240 780
rect -150 760 -90 810
rect 120 780 180 810
rect -1490 613 -1350 640
rect -1490 567 -1443 613
rect -1397 567 -1350 613
rect -1490 540 -1350 567
rect -1490 490 -1430 540
rect -1300 490 -1240 660
rect -870 490 -810 660
rect -730 580 -670 670
rect -560 610 -490 720
rect -340 697 -313 743
rect -267 697 -240 743
rect -340 660 -240 697
rect -170 718 -70 760
rect -170 672 -143 718
rect -97 672 -70 718
rect -170 630 -70 672
rect -20 728 70 760
rect -20 682 2 728
rect 48 682 70 728
rect -560 588 -430 610
rect -730 520 -620 580
rect -560 542 -538 588
rect -492 542 -430 588
rect -150 580 -90 630
rect -560 520 -430 542
rect -680 490 -620 520
rect -490 490 -430 520
rect -340 520 -90 580
rect -20 540 70 682
rect -340 490 -280 520
rect 10 490 70 540
rect 120 753 240 780
rect 120 707 157 753
rect 203 707 240 753
rect 120 680 240 707
rect 120 490 180 680
rect 310 490 370 810
rect 790 730 850 800
rect 1210 780 1270 810
rect 700 678 850 730
rect 700 632 752 678
rect 798 632 850 678
rect 1110 743 1270 780
rect 1110 697 1152 743
rect 1198 697 1270 743
rect 1110 660 1270 697
rect 1370 780 1430 810
rect 1370 748 1510 780
rect 1370 702 1432 748
rect 1478 702 1510 748
rect 1370 670 1510 702
rect 700 580 850 632
rect 790 490 850 580
rect 1180 490 1240 660
rect 1370 490 1430 670
rect 1560 650 1620 810
rect 1710 710 1770 810
rect 1900 760 1960 810
rect 2090 780 2150 810
rect 2090 753 2210 780
rect 1710 650 1960 710
rect 1560 618 1660 650
rect 1560 572 1587 618
rect 1633 572 1660 618
rect 1560 540 1660 572
rect 1900 630 1960 650
rect 2090 707 2127 753
rect 2173 707 2210 753
rect 2090 680 2210 707
rect 2280 700 2340 810
rect 2540 700 2660 730
rect 2280 693 2660 700
rect 1900 608 2020 630
rect 1900 562 1937 608
rect 1983 562 2020 608
rect 1900 540 2020 562
rect 1560 490 1620 540
rect 1710 490 1770 540
rect 1900 490 1960 540
rect 2090 490 2150 680
rect 2280 647 2577 693
rect 2623 647 2660 693
rect 2280 640 2660 647
rect 2280 490 2340 640
rect 2540 610 2660 640
rect -1490 270 -1430 320
rect -1300 270 -1240 320
rect -870 270 -810 320
rect -680 270 -620 320
rect -490 270 -430 320
rect -340 270 -280 320
rect 10 220 70 320
rect 120 270 180 320
rect 310 220 370 320
rect 790 270 850 320
rect 1180 270 1240 320
rect 1370 270 1430 320
rect 1560 270 1620 320
rect 1710 220 1770 320
rect 1900 270 1960 320
rect 2090 270 2150 320
rect 2280 220 2340 320
rect 10 160 2340 220
<< polycontact >>
rect -1073 687 -1027 733
rect -698 702 -652 748
rect -1443 567 -1397 613
rect -313 697 -267 743
rect -143 672 -97 718
rect 2 682 48 728
rect -538 542 -492 588
rect 157 707 203 753
rect 752 632 798 678
rect 1152 697 1198 743
rect 1432 702 1478 748
rect 1587 572 1633 618
rect 2127 707 2173 753
rect 1937 562 1983 608
rect 2577 647 2623 693
<< metal1 >>
rect -1690 1318 3840 1370
rect -1690 1272 -1543 1318
rect -1497 1272 2420 1318
rect 2560 1272 3840 1318
rect -1690 1268 3840 1272
rect -1690 1230 647 1268
rect -1590 1093 -1520 1150
rect -1590 1047 -1578 1093
rect -1532 1047 -1520 1093
rect -1590 750 -1520 1047
rect -1400 1093 -1329 1230
rect -1400 1047 -1388 1093
rect -1342 1047 -1329 1093
rect -1400 940 -1329 1047
rect -1210 1093 -1140 1150
rect -1210 1047 -1198 1093
rect -1152 1047 -1140 1093
rect -1400 913 -1330 940
rect -1400 867 -1388 913
rect -1342 867 -1330 913
rect -1400 810 -1330 867
rect -1210 913 -1140 1047
rect -1210 867 -1198 913
rect -1152 867 -1140 913
rect -1670 600 -1520 750
rect -1210 640 -1140 867
rect -1090 1093 -870 1150
rect -1090 1047 -928 1093
rect -882 1047 -870 1093
rect -1090 1020 -870 1047
rect -1090 733 -1010 1020
rect -1090 687 -1073 733
rect -1027 687 -1010 733
rect -1090 660 -1010 687
rect -940 913 -870 1020
rect -620 1093 -550 1230
rect -620 1047 -608 1093
rect -562 1047 -550 1093
rect -620 990 -550 1047
rect -500 1093 -180 1150
rect -500 1047 -248 1093
rect -202 1047 -180 1093
rect -500 990 -180 1047
rect 210 1093 280 1230
rect 600 1222 647 1230
rect 693 1250 3840 1268
rect 693 1230 2660 1250
rect 693 1222 760 1230
rect 600 1200 760 1222
rect 210 1047 222 1093
rect 268 1047 280 1093
rect 210 990 280 1047
rect 330 1020 640 1150
rect -500 940 -440 990
rect 330 940 400 1020
rect -940 867 -928 913
rect -882 867 -870 913
rect -1590 428 -1520 600
rect -1470 613 -1140 640
rect -1470 567 -1443 613
rect -1397 567 -1140 613
rect -1470 540 -1140 567
rect -940 610 -870 867
rect -730 880 -440 940
rect -730 748 -620 880
rect -730 702 -698 748
rect -652 720 -620 748
rect -340 820 70 940
rect -340 743 -240 820
rect -652 702 -390 720
rect -730 660 -390 702
rect -340 697 -313 743
rect -267 697 -240 743
rect -340 660 -240 697
rect -150 718 -70 760
rect -150 672 -143 718
rect -97 672 -70 718
rect -940 588 -490 610
rect -940 542 -538 588
rect -492 542 -490 588
rect -940 540 -490 542
rect -1590 382 -1578 428
rect -1532 382 -1520 428
rect -1590 320 -1520 382
rect -1400 428 -1329 494
rect -1400 382 -1388 428
rect -1342 382 -1329 428
rect -1400 240 -1329 382
rect -1210 428 -1140 540
rect -780 520 -490 540
rect -1210 382 -1198 428
rect -1152 382 -1140 428
rect -1210 320 -1140 382
rect -970 428 -900 490
rect -970 382 -958 428
rect -912 382 -900 428
rect -970 240 -900 382
rect -780 428 -700 520
rect -780 382 -768 428
rect -722 382 -700 428
rect -780 320 -700 382
rect -590 418 -520 470
rect -590 372 -578 418
rect -532 372 -520 418
rect -590 240 -520 372
rect -440 430 -390 660
rect -150 530 -70 672
rect 0 728 70 820
rect 0 682 2 728
rect 48 682 70 728
rect 120 880 400 940
rect 450 913 520 970
rect 120 753 240 880
rect 120 707 157 753
rect 203 707 240 753
rect 120 700 240 707
rect 450 867 462 913
rect 508 867 520 913
rect 570 940 640 1020
rect 690 1083 760 1200
rect 690 1037 702 1083
rect 748 1037 760 1083
rect 1100 1093 1350 1150
rect 1100 1080 1122 1093
rect 690 990 760 1037
rect 810 1047 1122 1080
rect 1168 1047 1350 1093
rect 810 1030 1350 1047
rect 810 1020 1180 1030
rect 810 940 870 1020
rect 570 870 870 940
rect 920 913 1060 970
rect 0 580 70 682
rect 450 530 520 867
rect 920 867 932 913
rect 978 867 1060 913
rect 920 810 1060 867
rect 1110 913 1180 1020
rect 1110 867 1122 913
rect 1168 867 1180 913
rect 1110 810 1180 867
rect 1000 760 1060 810
rect 1000 743 1240 760
rect 700 678 850 730
rect 700 632 752 678
rect 798 632 850 678
rect 700 580 850 632
rect 1000 697 1152 743
rect 1198 697 1240 743
rect 1000 680 1240 697
rect 1000 610 1060 680
rect -150 470 520 530
rect 920 540 1060 610
rect 1290 630 1350 1030
rect 1460 1093 1530 1230
rect 1460 1047 1472 1093
rect 1518 1047 1530 1093
rect 1460 913 1530 1047
rect 1460 867 1472 913
rect 1518 867 1530 913
rect 1460 810 1530 867
rect 1580 1093 1870 1150
rect 1580 1047 1812 1093
rect 1858 1047 1870 1093
rect 1580 1030 1870 1047
rect 1580 760 1650 1030
rect 1400 748 1650 760
rect 1400 702 1432 748
rect 1478 702 1650 748
rect 1400 680 1650 702
rect 1800 913 1870 1030
rect 1800 867 1812 913
rect 1858 867 1870 913
rect 1290 618 1660 630
rect 1290 572 1587 618
rect 1633 572 1660 618
rect 1290 540 1660 572
rect -440 408 -180 430
rect 400 428 520 470
rect -440 362 -248 408
rect -202 362 -180 408
rect -440 320 -180 362
rect 210 393 280 420
rect 210 347 222 393
rect 268 347 280 393
rect 210 240 280 347
rect 400 382 412 428
rect 458 382 520 428
rect 400 320 520 382
rect 690 428 760 490
rect 690 382 702 428
rect 748 382 760 428
rect 690 240 760 382
rect 920 428 990 540
rect 1290 490 1350 540
rect 920 382 932 428
rect 978 382 990 428
rect 920 320 990 382
rect 1080 428 1150 490
rect 1080 382 1092 428
rect 1138 382 1150 428
rect 1080 240 1150 382
rect 1270 428 1350 490
rect 1270 382 1282 428
rect 1328 382 1350 428
rect 1270 320 1350 382
rect 1460 428 1530 490
rect 1460 382 1472 428
rect 1518 382 1530 428
rect 1460 240 1530 382
rect 1800 428 1870 867
rect 2180 1093 2250 1230
rect 2180 1047 2192 1093
rect 2238 1047 2250 1093
rect 2180 913 2250 1047
rect 2180 867 2192 913
rect 2238 867 2250 913
rect 2180 810 2250 867
rect 2300 1020 2660 1150
rect 2300 760 2370 1020
rect 2090 753 2370 760
rect 2090 707 2127 753
rect 2173 707 2370 753
rect 2090 700 2370 707
rect 2420 913 2490 970
rect 2420 867 2432 913
rect 2478 867 2490 913
rect 2420 630 2490 867
rect 1920 608 2490 630
rect 2540 693 2660 730
rect 2540 647 2577 693
rect 2623 647 2660 693
rect 2540 610 2660 647
rect 1920 562 1937 608
rect 1983 562 2490 608
rect 1920 540 2490 562
rect 2420 490 2490 540
rect 2760 520 2880 610
rect 3140 520 3260 610
rect 3490 540 3640 630
rect 1800 382 1812 428
rect 1858 382 1870 428
rect 1800 320 1870 382
rect 2180 428 2250 490
rect 2180 382 2192 428
rect 2238 382 2250 428
rect 2180 240 2250 382
rect 2370 428 2490 490
rect 2370 382 2382 428
rect 2428 382 2490 428
rect 2370 320 2490 382
rect -1690 220 2660 240
rect -1690 198 3840 220
rect -1690 152 -1603 198
rect -1557 152 -830 198
rect -690 152 -220 198
rect -80 152 2420 198
rect 2560 152 3840 198
rect -1690 100 3840 152
use mux_as_component  mux_as_component_0
timestamp 1756740009
transform 1 0 2330 0 1 350
box 330 -250 1510 1020
<< labels >>
flabel metal1 s 2760 520 2880 610 0 FreeSans 600 0 0 0 A
port 3 nsew
flabel metal1 s 3140 520 3260 610 0 FreeSans 600 0 0 0 B
port 4 nsew
flabel metal1 s 3490 540 3640 630 0 FreeSans 600 0 0 0 S
port 5 nsew
flabel metal1 s 2540 610 2660 730 0 FreeSans 600 0 0 0 CLK
port 6 nsew
flabel metal1 s 700 580 850 730 0 FreeSans 600 0 0 0 RN
port 7 nsew
flabel metal1 s -1670 600 -1520 750 0 FreeSans 600 0 0 0 Q
port 8 nsew
flabel metal1 s -1690 100 3840 240 0 FreeSans 480 0 0 0 VSS
port 1 nsew
flabel metal1 s -1690 1230 3840 1370 0 FreeSans 480 0 0 0 VDD
port 0 nsew
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1756208311
<< nwell >>
rect 1308 188 1366 200
<< ndiffc >>
rect 1155 -195 1201 -51
<< polysilicon >>
rect 246 735 634 795
rect 246 675 306 735
rect 574 676 634 735
rect 246 140 306 267
rect 410 266 470 315
rect 410 247 510 266
rect 410 187 430 247
rect 490 187 510 247
rect 410 166 510 187
rect 246 122 351 140
rect 246 62 278 122
rect 338 62 351 122
rect 246 40 351 62
rect 246 -18 306 40
rect 410 -45 470 166
rect 738 113 798 269
rect 862 248 962 270
rect 862 188 884 248
rect 944 188 962 248
rect 862 170 962 188
rect 518 69 798 113
rect 518 9 532 69
rect 592 54 798 69
rect 592 9 634 54
rect 518 -14 634 9
rect 902 6 962 170
rect 1066 161 1126 255
rect 1013 139 1126 161
rect 1013 79 1036 139
rect 1096 79 1126 139
rect 1013 59 1126 79
rect 1066 0 1126 59
rect 1230 134 1290 255
rect 1230 114 1350 134
rect 1230 54 1269 114
rect 1329 54 1350 114
rect 1230 34 1350 54
rect 1230 -41 1290 34
rect 246 -312 306 -252
rect 738 -312 798 -252
rect 246 -372 798 -312
<< polycontact >>
rect 430 187 490 247
rect 278 62 338 122
rect 884 188 944 248
rect 532 9 592 69
rect 1036 79 1096 139
rect 1269 54 1329 114
<< metal1 >>
rect 0 706 1551 847
rect 96 61 110 121
rect 170 -182 218 544
rect 334 303 382 706
rect 410 187 430 247
rect 490 187 510 247
rect 662 139 710 544
rect 990 294 1038 706
rect 1318 248 1366 630
rect 862 188 884 248
rect 944 188 1366 248
rect 662 138 751 139
rect 264 62 278 122
rect 338 62 364 122
rect 662 80 677 138
rect 735 80 751 138
rect 662 79 751 80
rect 1007 79 1036 139
rect 1096 79 1107 139
rect 513 9 532 69
rect 592 9 615 69
rect 334 -282 382 -41
rect 662 -182 710 79
rect 990 -282 1038 -42
rect 1155 -51 1201 188
rect 1248 54 1269 114
rect 1329 54 1348 114
rect 1155 -206 1201 -195
rect 1318 -282 1366 -28
rect 0 -423 1551 -282
<< via1 >>
rect 110 61 170 121
rect 677 80 735 138
<< metal2 >>
rect 410 178 510 258
rect 677 142 735 150
rect 675 139 737 142
rect 1024 139 1126 149
rect 671 138 1126 139
rect 99 121 179 132
rect 99 61 110 121
rect 170 61 179 121
rect 99 52 179 61
rect 264 53 364 133
rect 671 80 677 138
rect 735 80 1126 138
rect 110 -81 170 52
rect 513 0 614 80
rect 671 79 1126 80
rect 675 77 737 79
rect 677 68 735 77
rect 1024 69 1126 79
rect 1237 45 1349 124
rect 533 -81 593 0
rect 110 -141 593 -81
use nfet_03v3_CWXVHP  nfet_03v3_CWXVHP_0
timestamp 1756208265
transform 1 0 768 0 1 -123
box -610 -129 610 129
use pfet_03v3_XSU2S3  pfet_03v3_XSU2S3_0
timestamp 1756208265
transform 1 0 768 0 1 462
box -696 -300 696 300
<< end >>

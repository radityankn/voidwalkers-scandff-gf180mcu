magic
tech gf180mcuD
magscale 1 5
timestamp 1756545041
<< error_p >>
rect -25 575 30 685
rect -73 405 30 575
rect -40 335 -30 338
rect -48 315 -30 335
rect -25 325 30 405
rect -25 270 -7 315
rect -30 160 -2 245
rect -49 110 -45 134
rect -25 80 -6 110
rect -25 50 -7 80
<< nwell >>
rect -745 325 -30 685
rect -25 325 1305 685
<< pwell >>
rect -745 50 -30 325
rect -25 270 1305 325
rect -25 260 980 270
rect 1045 260 1075 270
rect 1140 260 1170 270
rect 1210 260 1305 270
rect -25 50 1305 260
<< nmos >>
rect -630 160 -600 245
rect -435 160 -405 245
rect -340 160 -310 245
rect -245 160 -215 245
rect -170 160 -140 245
rect -75 160 -45 245
rect 20 160 50 245
rect 115 160 145 245
rect 395 160 425 245
rect 590 160 620 245
rect 685 160 715 245
rect 780 160 810 245
rect 855 160 885 245
rect 950 160 980 245
rect 1045 160 1075 245
rect 1140 160 1170 245
<< pmos >>
rect -630 405 -600 575
rect -420 405 -390 575
rect -340 405 -310 575
rect -245 405 -215 575
rect -170 405 -140 575
rect -75 405 -45 575
rect 20 405 50 575
rect 115 405 145 575
rect 395 405 425 575
rect 605 405 635 575
rect 685 405 715 575
rect 780 405 810 575
rect 855 405 885 575
rect 950 405 980 575
rect 1045 405 1075 575
rect 1140 405 1170 575
<< ndiff >>
rect -685 235 -630 245
rect -685 170 -675 235
rect -650 170 -630 235
rect -685 160 -630 170
rect -600 235 -525 245
rect -600 170 -560 235
rect -535 170 -525 235
rect -600 160 -525 170
rect -490 235 -435 245
rect -490 170 -480 235
rect -455 170 -435 235
rect -490 160 -435 170
rect -405 235 -340 245
rect -405 170 -390 235
rect -355 170 -340 235
rect -405 160 -340 170
rect -310 235 -245 245
rect -310 170 -290 235
rect -265 170 -245 235
rect -310 160 -245 170
rect -215 160 -170 245
rect -140 235 -75 245
rect -140 170 -120 235
rect -95 170 -75 235
rect -140 160 -75 170
rect -45 160 -30 245
rect -25 160 20 245
rect 50 235 115 245
rect 50 170 70 235
rect 95 170 115 235
rect 50 160 115 170
rect 145 235 235 245
rect 145 170 165 235
rect 190 170 235 235
rect 145 160 235 170
rect 340 235 395 245
rect 340 170 350 235
rect 375 170 395 235
rect 340 160 395 170
rect 425 235 500 245
rect 425 170 465 235
rect 490 170 500 235
rect 425 160 500 170
rect 535 235 590 245
rect 535 170 545 235
rect 570 170 590 235
rect 535 160 590 170
rect 620 235 685 245
rect 620 170 635 235
rect 670 170 685 235
rect 620 160 685 170
rect 715 235 780 245
rect 715 170 735 235
rect 760 170 780 235
rect 715 160 780 170
rect 810 160 855 245
rect 885 235 950 245
rect 885 170 905 235
rect 930 170 950 235
rect 885 160 950 170
rect 980 160 1045 245
rect 1075 235 1140 245
rect 1075 170 1095 235
rect 1120 170 1140 235
rect 1075 160 1140 170
rect 1170 235 1260 245
rect 1170 170 1190 235
rect 1215 170 1260 235
rect 1170 160 1260 170
<< pdiff >>
rect -685 565 -630 575
rect -685 505 -675 565
rect -650 505 -630 565
rect -685 475 -630 505
rect -685 415 -675 475
rect -650 415 -630 475
rect -685 405 -630 415
rect -600 475 -525 575
rect -600 415 -560 475
rect -535 415 -525 475
rect -600 405 -525 415
rect -475 565 -420 575
rect -475 505 -465 565
rect -440 505 -420 565
rect -475 475 -420 505
rect -475 415 -465 475
rect -440 415 -420 475
rect -475 405 -420 415
rect -390 405 -340 575
rect -310 565 -245 575
rect -310 505 -290 565
rect -265 505 -245 565
rect -310 475 -245 505
rect -310 415 -290 475
rect -265 415 -245 475
rect -310 405 -245 415
rect -215 405 -170 575
rect -140 565 -75 575
rect -140 505 -120 565
rect -95 505 -75 565
rect -140 475 -75 505
rect -140 415 -120 475
rect -95 415 -75 475
rect -140 405 -75 415
rect -45 405 -30 575
rect -25 405 20 575
rect 50 565 115 575
rect 50 505 70 565
rect 95 505 115 565
rect 50 475 115 505
rect 50 415 70 475
rect 95 415 115 475
rect 50 405 115 415
rect 145 475 235 575
rect 145 415 190 475
rect 215 415 235 475
rect 145 405 235 415
rect 340 565 395 575
rect 340 505 350 565
rect 375 505 395 565
rect 340 405 395 505
rect 425 475 500 575
rect 425 415 465 475
rect 490 415 500 475
rect 425 405 500 415
rect 550 565 605 575
rect 550 505 560 565
rect 585 505 605 565
rect 550 475 605 505
rect 550 415 560 475
rect 585 415 605 475
rect 550 405 605 415
rect 635 405 685 575
rect 715 565 780 575
rect 715 505 735 565
rect 760 505 780 565
rect 715 475 780 505
rect 715 415 735 475
rect 760 415 780 475
rect 715 405 780 415
rect 810 405 855 575
rect 885 565 950 575
rect 885 505 905 565
rect 930 505 950 565
rect 885 475 950 505
rect 885 415 905 475
rect 930 415 950 475
rect 885 405 950 415
rect 980 405 1045 575
rect 1075 565 1140 575
rect 1075 505 1095 565
rect 1120 505 1140 565
rect 1075 475 1140 505
rect 1075 415 1095 475
rect 1120 415 1140 475
rect 1075 405 1140 415
rect 1170 475 1260 575
rect 1170 415 1215 475
rect 1240 415 1260 475
rect 1170 405 1260 415
<< ndiffc >>
rect -675 170 -650 235
rect -560 170 -535 235
rect -480 170 -455 235
rect -390 170 -355 235
rect -290 170 -265 235
rect -120 170 -95 235
rect 70 170 95 235
rect 165 170 190 235
rect 350 170 375 235
rect 465 170 490 235
rect 545 170 570 235
rect 635 170 670 235
rect 735 170 760 235
rect 905 170 930 235
rect 1095 170 1120 235
rect 1190 170 1215 235
<< pdiffc >>
rect -675 505 -650 565
rect -675 415 -650 475
rect -560 415 -535 475
rect -465 505 -440 565
rect -465 415 -440 475
rect -290 505 -265 565
rect -290 415 -265 475
rect -120 505 -95 565
rect -120 415 -95 475
rect 70 505 95 565
rect 70 415 95 475
rect 190 415 215 475
rect 350 505 375 565
rect 465 415 490 475
rect 560 505 585 565
rect 560 415 585 475
rect 735 505 760 565
rect 735 415 760 475
rect 905 505 930 565
rect 905 415 930 475
rect 1095 505 1120 565
rect 1095 415 1120 475
rect 1215 415 1240 475
<< polysilicon >>
rect -170 625 -30 655
rect -25 625 145 655
rect -630 575 -600 600
rect -420 575 -390 600
rect -340 575 -310 600
rect -245 575 -215 600
rect -170 575 -140 625
rect -75 575 -45 600
rect 20 575 50 600
rect 115 575 145 625
rect 950 625 1170 655
rect 395 575 425 600
rect 605 575 635 600
rect 685 575 715 600
rect 780 575 810 600
rect 855 575 885 600
rect 950 575 980 625
rect 1045 575 1075 600
rect 1140 575 1170 625
rect -630 245 -600 405
rect -420 390 -390 405
rect -470 380 -390 390
rect -470 340 -460 380
rect -415 340 -390 380
rect -470 330 -390 340
rect -340 390 -310 405
rect -340 380 -270 390
rect -340 345 -315 380
rect -280 345 -270 380
rect -340 335 -270 345
rect -435 245 -405 330
rect -340 245 -310 335
rect -245 325 -215 405
rect -170 380 -140 405
rect -75 390 -45 405
rect 20 390 50 405
rect -75 380 -30 390
rect -75 335 -65 380
rect -40 335 -30 380
rect -75 325 -30 335
rect 20 380 80 390
rect 20 350 30 380
rect 70 350 80 380
rect 20 340 80 350
rect -245 315 -195 325
rect -245 280 -235 315
rect -205 280 -195 315
rect -245 270 -195 280
rect -170 295 -45 325
rect -245 245 -215 270
rect -170 245 -140 295
rect -75 245 -45 270
rect 20 245 50 340
rect 115 245 145 405
rect 395 245 425 405
rect 605 390 635 405
rect 555 380 635 390
rect 555 340 565 380
rect 610 340 635 380
rect 555 330 635 340
rect 685 390 715 405
rect 685 380 755 390
rect 685 345 710 380
rect 745 345 755 380
rect 685 335 755 345
rect 590 245 620 330
rect 685 245 715 335
rect 780 325 810 405
rect 855 355 885 405
rect 950 380 980 405
rect 1045 390 1075 405
rect 1045 380 1105 390
rect 855 325 980 355
rect 780 315 830 325
rect 780 280 790 315
rect 820 280 830 315
rect 780 270 830 280
rect 950 315 980 325
rect 1045 350 1055 380
rect 1095 350 1105 380
rect 1045 340 1105 350
rect 1140 350 1170 405
rect 950 305 1010 315
rect 950 280 960 305
rect 1000 280 1010 305
rect 950 270 1010 280
rect 780 245 810 270
rect 855 245 885 270
rect 950 245 980 270
rect 1045 245 1075 340
rect 1140 320 1290 350
rect 1140 245 1170 320
rect -630 135 -600 160
rect -435 135 -405 160
rect -340 135 -310 160
rect -245 135 -215 160
rect -170 135 -140 160
rect -75 110 -45 160
rect 20 135 50 160
rect 115 110 145 160
rect 395 135 425 160
rect 590 135 620 160
rect 685 135 715 160
rect 780 135 810 160
rect 855 110 885 160
rect 950 135 980 160
rect 1045 135 1075 160
rect 1140 110 1170 160
rect -75 80 -30 110
rect -25 80 1170 110
<< polycontact >>
rect -460 340 -415 380
rect -315 345 -280 380
rect -65 335 -40 380
rect 30 350 70 380
rect -235 280 -205 315
rect 565 340 610 380
rect 710 345 745 380
rect 790 280 820 315
rect 1055 350 1095 380
rect 960 280 1000 305
<< metal1 >>
rect -745 625 -30 685
rect -25 625 1305 685
rect -680 565 -645 625
rect -680 505 -675 565
rect -650 505 -645 565
rect -680 475 -645 505
rect -680 415 -675 475
rect -650 415 -645 475
rect -680 405 -645 415
rect -620 565 -350 575
rect -620 510 -465 565
rect -620 300 -590 510
rect -470 505 -465 510
rect -440 515 -350 565
rect -440 505 -435 515
rect -565 475 -495 485
rect -565 415 -560 475
rect -535 415 -495 475
rect -565 405 -495 415
rect -470 475 -435 505
rect -470 415 -465 475
rect -440 415 -435 475
rect -470 405 -435 415
rect -525 380 -495 405
rect -525 340 -460 380
rect -415 340 -405 380
rect -525 305 -495 340
rect -745 270 -590 300
rect -565 270 -495 305
rect -380 315 -350 515
rect -295 565 -260 625
rect -295 505 -290 565
rect -265 505 -260 565
rect -295 475 -260 505
rect -295 415 -290 475
rect -265 415 -260 475
rect -295 405 -260 415
rect -235 565 -90 575
rect -235 515 -120 565
rect -235 380 -200 515
rect -325 345 -315 380
rect -280 345 -200 380
rect -325 340 -200 345
rect -125 505 -120 515
rect -95 505 -90 565
rect -125 475 -90 505
rect -125 415 -120 475
rect -95 415 -90 475
rect -380 280 -235 315
rect -205 280 -195 315
rect -380 270 -195 280
rect -680 235 -645 245
rect -680 170 -675 235
rect -650 170 -645 235
rect -680 110 -645 170
rect -565 235 -530 270
rect -380 245 -350 270
rect -565 170 -560 235
rect -535 170 -530 235
rect -565 160 -530 170
rect -485 235 -450 245
rect -485 170 -480 235
rect -455 170 -450 235
rect -485 110 -450 170
rect -390 235 -350 245
rect -355 170 -350 235
rect -390 160 -350 170
rect -295 235 -260 245
rect -295 170 -290 235
rect -265 170 -260 235
rect -295 110 -260 170
rect -125 235 -90 415
rect 65 565 100 625
rect 65 505 70 565
rect 95 505 100 565
rect 65 475 100 505
rect 65 415 70 475
rect 95 415 100 475
rect 65 405 100 415
rect 125 510 280 575
rect -65 380 -30 390
rect 125 380 160 510
rect -40 335 -30 380
rect 20 350 30 380
rect 70 350 160 380
rect 185 475 220 485
rect 185 415 190 475
rect 215 415 220 475
rect 245 470 280 510
rect 345 565 380 625
rect 345 505 350 565
rect 375 505 380 565
rect 345 495 380 505
rect 405 565 675 575
rect 405 510 560 565
rect 405 470 435 510
rect 555 505 560 510
rect 585 515 675 565
rect 585 505 590 515
rect 245 435 435 470
rect -65 270 -30 335
rect 185 315 220 415
rect -25 270 220 315
rect 405 300 435 435
rect 460 475 530 485
rect 460 415 465 475
rect 490 415 530 475
rect 460 405 530 415
rect 555 475 590 505
rect 555 415 560 475
rect 585 415 590 475
rect 555 405 590 415
rect 500 380 530 405
rect 500 340 565 380
rect 610 340 620 380
rect 500 305 530 340
rect 280 270 435 300
rect 460 270 530 305
rect 645 315 675 515
rect 730 565 765 625
rect 730 505 735 565
rect 760 505 765 565
rect 730 475 765 505
rect 730 415 735 475
rect 760 415 765 475
rect 730 405 765 415
rect 790 565 935 575
rect 790 515 905 565
rect 790 380 825 515
rect 700 345 710 380
rect 745 345 825 380
rect 700 340 825 345
rect 900 505 905 515
rect 930 505 935 565
rect 900 475 935 505
rect 900 415 905 475
rect 930 415 935 475
rect 645 280 790 315
rect 820 280 830 315
rect 645 270 830 280
rect 185 245 220 270
rect -125 170 -120 235
rect -95 170 -90 235
rect -125 160 -90 170
rect 65 235 100 245
rect 65 170 70 235
rect 95 170 100 235
rect -75 110 -45 140
rect 65 110 100 170
rect 160 235 220 245
rect 160 170 165 235
rect 190 170 220 235
rect 160 160 220 170
rect 345 235 380 245
rect 345 170 350 235
rect 375 170 380 235
rect 345 110 380 170
rect 460 235 495 270
rect 645 245 675 270
rect 460 170 465 235
rect 490 170 495 235
rect 460 160 495 170
rect 540 235 575 245
rect 540 170 545 235
rect 570 170 575 235
rect 540 110 575 170
rect 635 235 675 245
rect 670 170 675 235
rect 635 160 675 170
rect 730 235 765 245
rect 730 170 735 235
rect 760 170 765 235
rect 730 110 765 170
rect 900 235 935 415
rect 1090 565 1125 625
rect 1090 505 1095 565
rect 1120 505 1125 565
rect 1090 475 1125 505
rect 1090 415 1095 475
rect 1120 415 1125 475
rect 1090 405 1125 415
rect 1150 510 1260 575
rect 1150 380 1185 510
rect 1045 350 1055 380
rect 1095 350 1185 380
rect 1210 475 1245 485
rect 1210 415 1215 475
rect 1240 415 1245 475
rect 1210 315 1245 415
rect 960 305 1245 315
rect 1000 280 1245 305
rect 960 270 1245 280
rect 1210 245 1245 270
rect 900 170 905 235
rect 930 170 935 235
rect 900 160 935 170
rect 1090 235 1125 245
rect 1090 170 1095 235
rect 1120 170 1125 235
rect 1090 110 1125 170
rect 1185 235 1245 245
rect 1185 170 1190 235
rect 1215 170 1245 235
rect 1185 160 1245 170
rect -745 50 -30 110
rect -25 50 1305 110
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1756212155
<< nmos >>
rect -112 -85 -52 85
rect 52 -85 112 85
<< ndiff >>
rect -200 72 -112 85
rect -200 -72 -187 72
rect -141 -72 -112 72
rect -200 -85 -112 -72
rect -52 72 52 85
rect -52 -72 -23 72
rect 23 -72 52 72
rect -52 -85 52 -72
rect 112 72 200 85
rect 112 -72 141 72
rect 187 -72 200 72
rect 112 -85 200 -72
<< ndiffc >>
rect -187 -72 -141 72
rect -23 -72 23 72
rect 141 -72 187 72
<< polysilicon >>
rect -112 85 -52 129
rect 52 85 112 129
rect -112 -129 -52 -85
rect 52 -129 112 -85
<< metal1 >>
rect -187 72 -141 83
rect -187 -83 -141 -72
rect -23 72 23 83
rect -23 -83 23 -72
rect 141 72 187 83
rect 141 -83 187 -72
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.85 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1756212155
<< nwell >>
rect -204 -300 204 300
<< pmos >>
rect -30 -170 30 170
<< pdiff >>
rect -118 157 -30 170
rect -118 -157 -105 157
rect -59 -157 -30 157
rect -118 -170 -30 -157
rect 30 157 118 170
rect 30 -157 59 157
rect 105 -157 118 157
rect 30 -170 118 -157
<< pdiffc >>
rect -105 -157 -59 157
rect 59 -157 105 157
<< polysilicon >>
rect -30 170 30 214
rect -30 -214 30 -170
<< metal1 >>
rect -105 157 -59 168
rect -105 -168 -59 -157
rect 59 157 105 168
rect 59 -168 105 -157
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.7 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>

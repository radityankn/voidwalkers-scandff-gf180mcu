magic
tech gf180mcuD
magscale 1 10
timestamp 1756235029
<< nwell >>
rect -614 -300 614 300
<< pmos >>
rect -440 -170 -380 170
rect -276 -170 -216 170
rect -112 -170 -52 170
rect 52 -170 112 170
rect 216 -170 276 170
rect 380 -170 440 170
<< pdiff >>
rect -528 157 -440 170
rect -528 -157 -515 157
rect -469 -157 -440 157
rect -528 -170 -440 -157
rect -380 -170 -276 170
rect -216 157 -112 170
rect -216 -157 -187 157
rect -141 -157 -112 157
rect -216 -170 -112 -157
rect -52 -170 52 170
rect 112 157 216 170
rect 112 -157 141 157
rect 187 -157 216 157
rect 112 -170 216 -157
rect 276 -170 380 170
rect 440 157 528 170
rect 440 -157 469 157
rect 515 -157 528 157
rect 440 -170 528 -157
<< pdiffc >>
rect -515 -157 -469 157
rect -187 -157 -141 157
rect 141 -157 187 157
rect 469 -157 515 157
<< polysilicon >>
rect -440 170 -380 214
rect -276 170 -216 214
rect -112 170 -52 214
rect 52 170 112 214
rect 216 170 276 214
rect 380 170 440 214
rect -440 -214 -380 -170
rect -276 -214 -216 -170
rect -112 -214 -52 -170
rect 52 -214 112 -170
rect 216 -214 276 -170
rect 380 -214 440 -170
<< metal1 >>
rect -515 157 -469 168
rect -515 -168 -469 -157
rect -187 157 -141 168
rect -187 -168 -141 -157
rect 141 157 187 168
rect 141 -168 187 -157
rect 469 157 515 168
rect 469 -168 515 -157
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.7 l 0.3 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1755195943
<< nwell >>
rect -1516 -300 1516 300
<< pmos >>
rect -1342 -170 -1282 170
rect -1178 -170 -1118 170
rect -1014 -170 -954 170
rect -850 -170 -790 170
rect -686 -170 -626 170
rect -522 -170 -462 170
rect -358 -170 -298 170
rect -194 -170 -134 170
rect -30 -170 30 170
rect 134 -170 194 170
rect 298 -170 358 170
rect 462 -170 522 170
rect 626 -170 686 170
rect 790 -170 850 170
rect 954 -170 1014 170
rect 1118 -170 1178 170
rect 1282 -170 1342 170
<< pdiff >>
rect -1430 157 -1342 170
rect -1430 -157 -1417 157
rect -1371 -157 -1342 157
rect -1430 -170 -1342 -157
rect -1282 157 -1178 170
rect -1282 -157 -1253 157
rect -1207 -157 -1178 157
rect -1282 -170 -1178 -157
rect -1118 157 -1014 170
rect -1118 -157 -1089 157
rect -1043 -157 -1014 157
rect -1118 -170 -1014 -157
rect -954 157 -850 170
rect -954 -157 -925 157
rect -879 -157 -850 157
rect -954 -170 -850 -157
rect -790 157 -686 170
rect -790 -157 -761 157
rect -715 -157 -686 157
rect -790 -170 -686 -157
rect -626 157 -522 170
rect -626 -157 -597 157
rect -551 -157 -522 157
rect -626 -170 -522 -157
rect -462 157 -358 170
rect -462 -157 -433 157
rect -387 -157 -358 157
rect -462 -170 -358 -157
rect -298 157 -194 170
rect -298 -157 -269 157
rect -223 -157 -194 157
rect -298 -170 -194 -157
rect -134 157 -30 170
rect -134 -157 -105 157
rect -59 -157 -30 157
rect -134 -170 -30 -157
rect 30 157 134 170
rect 30 -157 59 157
rect 105 -157 134 157
rect 30 -170 134 -157
rect 194 157 298 170
rect 194 -157 223 157
rect 269 -157 298 157
rect 194 -170 298 -157
rect 358 157 462 170
rect 358 -157 387 157
rect 433 -157 462 157
rect 358 -170 462 -157
rect 522 157 626 170
rect 522 -157 551 157
rect 597 -157 626 157
rect 522 -170 626 -157
rect 686 157 790 170
rect 686 -157 715 157
rect 761 -157 790 157
rect 686 -170 790 -157
rect 850 157 954 170
rect 850 -157 879 157
rect 925 -157 954 157
rect 850 -170 954 -157
rect 1014 157 1118 170
rect 1014 -157 1043 157
rect 1089 -157 1118 157
rect 1014 -170 1118 -157
rect 1178 157 1282 170
rect 1178 -157 1207 157
rect 1253 -157 1282 157
rect 1178 -170 1282 -157
rect 1342 157 1430 170
rect 1342 -157 1371 157
rect 1417 -157 1430 157
rect 1342 -170 1430 -157
<< pdiffc >>
rect -1417 -157 -1371 157
rect -1253 -157 -1207 157
rect -1089 -157 -1043 157
rect -925 -157 -879 157
rect -761 -157 -715 157
rect -597 -157 -551 157
rect -433 -157 -387 157
rect -269 -157 -223 157
rect -105 -157 -59 157
rect 59 -157 105 157
rect 223 -157 269 157
rect 387 -157 433 157
rect 551 -157 597 157
rect 715 -157 761 157
rect 879 -157 925 157
rect 1043 -157 1089 157
rect 1207 -157 1253 157
rect 1371 -157 1417 157
<< polysilicon >>
rect -1342 170 -1282 214
rect -1178 170 -1118 214
rect -1014 170 -954 214
rect -850 170 -790 214
rect -686 170 -626 214
rect -522 170 -462 214
rect -358 170 -298 214
rect -194 170 -134 214
rect -30 170 30 214
rect 134 170 194 214
rect 298 170 358 214
rect 462 170 522 214
rect 626 170 686 214
rect 790 170 850 214
rect 954 170 1014 214
rect 1118 170 1178 214
rect 1282 170 1342 214
rect -1342 -214 -1282 -170
rect -1178 -214 -1118 -170
rect -1014 -214 -954 -170
rect -850 -214 -790 -170
rect -686 -214 -626 -170
rect -522 -214 -462 -170
rect -358 -214 -298 -170
rect -194 -214 -134 -170
rect -30 -214 30 -170
rect 134 -214 194 -170
rect 298 -214 358 -170
rect 462 -214 522 -170
rect 626 -214 686 -170
rect 790 -214 850 -170
rect 954 -214 1014 -170
rect 1118 -214 1178 -170
rect 1282 -214 1342 -170
<< metal1 >>
rect -1417 157 -1371 168
rect -1417 -168 -1371 -157
rect -1253 157 -1207 168
rect -1253 -168 -1207 -157
rect -1089 157 -1043 168
rect -1089 -168 -1043 -157
rect -925 157 -879 168
rect -925 -168 -879 -157
rect -761 157 -715 168
rect -761 -168 -715 -157
rect -597 157 -551 168
rect -597 -168 -551 -157
rect -433 157 -387 168
rect -433 -168 -387 -157
rect -269 157 -223 168
rect -269 -168 -223 -157
rect -105 157 -59 168
rect -105 -168 -59 -157
rect 59 157 105 168
rect 59 -168 105 -157
rect 223 157 269 168
rect 223 -168 269 -157
rect 387 157 433 168
rect 387 -168 433 -157
rect 551 157 597 168
rect 551 -168 597 -157
rect 715 157 761 168
rect 715 -168 761 -157
rect 879 157 925 168
rect 879 -168 925 -157
rect 1043 157 1089 168
rect 1043 -168 1089 -157
rect 1207 157 1253 168
rect 1207 -168 1253 -157
rect 1371 157 1417 168
rect 1371 -168 1417 -157
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.7 l 0.3 m 1 nf 17 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1756675332
<< nwell >>
rect 330 300 1510 1020
<< pwell >>
rect 330 -250 1510 300
<< nmos >>
rect 580 -30 640 140
rect 770 -30 830 140
rect 1250 -30 1310 140
<< pmos >>
rect 580 460 640 800
rect 770 460 830 800
rect 1250 460 1310 800
<< ndiff >>
rect 459 120 580 140
rect 459 -10 490 120
rect 540 -10 580 120
rect 459 -30 580 -10
rect 640 120 770 140
rect 640 -10 680 120
rect 730 -10 770 120
rect 640 -30 770 -10
rect 830 120 960 140
rect 830 -10 870 120
rect 920 -10 960 120
rect 1120 120 1250 140
rect 830 -30 960 -10
rect 1120 -10 1160 120
rect 1210 -10 1250 120
rect 1120 -30 1250 -10
rect 1310 120 1420 140
rect 1310 -10 1350 120
rect 1400 -10 1420 120
rect 1310 -30 1420 -10
<< pdiff >>
rect 459 600 580 800
rect 459 480 490 600
rect 540 480 580 600
rect 459 460 580 480
rect 640 780 770 800
rect 640 660 680 780
rect 730 660 770 780
rect 640 600 770 660
rect 640 480 680 600
rect 730 480 770 600
rect 640 460 770 480
rect 830 780 960 800
rect 830 660 870 780
rect 920 660 960 780
rect 1120 780 1250 800
rect 830 600 960 660
rect 830 480 870 600
rect 920 480 960 600
rect 830 460 960 480
rect 1120 660 1160 780
rect 1210 660 1250 780
rect 1120 600 1250 660
rect 1120 480 1160 600
rect 1210 480 1250 600
rect 1120 460 1250 480
rect 1310 780 1420 800
rect 1310 660 1350 780
rect 1400 660 1420 780
rect 1310 600 1420 660
rect 1310 480 1350 600
rect 1400 480 1420 600
rect 1310 460 1420 480
<< ndiffc >>
rect 490 -10 540 120
rect 680 -10 730 120
rect 870 -10 920 120
rect 1160 -10 1210 120
rect 1350 -10 1400 120
<< pdiffc >>
rect 490 480 540 600
rect 680 660 730 780
rect 680 480 730 600
rect 870 660 920 780
rect 870 480 920 600
rect 1160 660 1210 780
rect 1160 480 1210 600
rect 1350 660 1400 780
rect 1350 480 1400 600
<< polysilicon >>
rect 770 850 1100 900
rect 580 800 640 850
rect 770 800 830 850
rect 1020 830 1100 850
rect 1020 719 1036 830
rect 1085 719 1100 830
rect 1250 800 1310 850
rect 1020 700 1100 719
rect 580 360 640 460
rect 770 410 830 460
rect 580 300 830 360
rect 770 290 830 300
rect 1250 290 1310 460
rect 770 270 1310 290
rect 770 210 1180 270
rect 1290 210 1310 270
rect 770 190 1310 210
rect 580 140 640 190
rect 770 140 830 190
rect 1250 140 1310 190
rect 1020 50 1100 70
rect 580 -130 640 -30
rect 770 -80 830 -30
rect 1020 -61 1036 50
rect 1085 -61 1100 50
rect 1020 -130 1100 -61
rect 1250 -80 1310 -30
rect 580 -190 1100 -130
<< polycontact >>
rect 1036 719 1085 830
rect 1180 210 1290 270
rect 1036 -61 1085 50
<< metal1 >>
rect 330 900 1510 1020
rect 1020 830 1100 850
rect 330 780 740 800
rect 330 670 680 780
rect 670 660 680 670
rect 730 660 740 780
rect 480 600 550 620
rect 480 480 490 600
rect 540 480 550 600
rect 480 260 550 480
rect 430 170 550 260
rect 480 120 550 170
rect 480 -10 490 120
rect 540 -10 550 120
rect 480 -30 550 -10
rect 670 600 740 660
rect 670 480 680 600
rect 730 480 740 600
rect 670 120 740 480
rect 860 780 930 800
rect 860 660 870 780
rect 920 660 930 780
rect 860 600 930 660
rect 860 480 870 600
rect 920 480 930 600
rect 860 260 930 480
rect 810 170 930 260
rect 670 -10 680 120
rect 730 -10 740 120
rect 670 -30 740 -10
rect 860 120 930 170
rect 860 -10 870 120
rect 920 -10 930 120
rect 860 -30 930 -10
rect 1020 719 1036 830
rect 1085 719 1100 830
rect 1020 410 1100 719
rect 1150 780 1220 900
rect 1150 660 1160 780
rect 1210 660 1220 780
rect 1150 600 1220 660
rect 1150 480 1160 600
rect 1210 480 1220 600
rect 1150 460 1220 480
rect 1340 780 1450 800
rect 1340 660 1350 780
rect 1400 660 1450 780
rect 1340 600 1450 660
rect 1340 480 1350 600
rect 1400 480 1450 600
rect 1340 460 1450 480
rect 1390 410 1450 460
rect 1020 330 1450 410
rect 1020 50 1100 330
rect 1160 270 1310 280
rect 1160 210 1180 270
rect 1290 210 1310 270
rect 1160 190 1310 210
rect 1390 140 1450 330
rect 1020 -61 1036 50
rect 1085 -61 1100 50
rect 1020 -80 1100 -61
rect 1150 120 1220 140
rect 1150 -10 1160 120
rect 1210 -10 1220 120
rect 1150 -130 1220 -10
rect 1340 120 1450 140
rect 1340 -10 1350 120
rect 1400 -10 1450 120
rect 1340 -30 1450 -10
rect 330 -250 1510 -130
<< end >>

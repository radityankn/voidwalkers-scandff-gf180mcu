magic
tech gf180mcuD
magscale 1 10
timestamp 1755195943
<< nwell >>
rect -2620 -300 2620 300
<< pmos >>
rect -2446 -170 -2386 170
rect -2144 -170 -2084 170
rect -1842 -170 -1782 170
rect -1540 -170 -1480 170
rect -1238 -170 -1178 170
rect -936 -170 -876 170
rect -634 -170 -574 170
rect -332 -170 -272 170
rect -30 -170 30 170
rect 272 -170 332 170
rect 574 -170 634 170
rect 876 -170 936 170
rect 1178 -170 1238 170
rect 1480 -170 1540 170
rect 1782 -170 1842 170
rect 2084 -170 2144 170
rect 2386 -170 2446 170
<< pdiff >>
rect -2534 157 -2446 170
rect -2534 -157 -2521 157
rect -2475 -157 -2446 157
rect -2534 -170 -2446 -157
rect -2386 157 -2298 170
rect -2386 -157 -2357 157
rect -2311 -157 -2298 157
rect -2386 -170 -2298 -157
rect -2232 157 -2144 170
rect -2232 -157 -2219 157
rect -2173 -157 -2144 157
rect -2232 -170 -2144 -157
rect -2084 157 -1996 170
rect -2084 -157 -2055 157
rect -2009 -157 -1996 157
rect -2084 -170 -1996 -157
rect -1930 157 -1842 170
rect -1930 -157 -1917 157
rect -1871 -157 -1842 157
rect -1930 -170 -1842 -157
rect -1782 157 -1694 170
rect -1782 -157 -1753 157
rect -1707 -157 -1694 157
rect -1782 -170 -1694 -157
rect -1628 157 -1540 170
rect -1628 -157 -1615 157
rect -1569 -157 -1540 157
rect -1628 -170 -1540 -157
rect -1480 157 -1392 170
rect -1480 -157 -1451 157
rect -1405 -157 -1392 157
rect -1480 -170 -1392 -157
rect -1326 157 -1238 170
rect -1326 -157 -1313 157
rect -1267 -157 -1238 157
rect -1326 -170 -1238 -157
rect -1178 157 -1090 170
rect -1178 -157 -1149 157
rect -1103 -157 -1090 157
rect -1178 -170 -1090 -157
rect -1024 157 -936 170
rect -1024 -157 -1011 157
rect -965 -157 -936 157
rect -1024 -170 -936 -157
rect -876 157 -788 170
rect -876 -157 -847 157
rect -801 -157 -788 157
rect -876 -170 -788 -157
rect -722 157 -634 170
rect -722 -157 -709 157
rect -663 -157 -634 157
rect -722 -170 -634 -157
rect -574 157 -486 170
rect -574 -157 -545 157
rect -499 -157 -486 157
rect -574 -170 -486 -157
rect -420 157 -332 170
rect -420 -157 -407 157
rect -361 -157 -332 157
rect -420 -170 -332 -157
rect -272 157 -184 170
rect -272 -157 -243 157
rect -197 -157 -184 157
rect -272 -170 -184 -157
rect -118 157 -30 170
rect -118 -157 -105 157
rect -59 -157 -30 157
rect -118 -170 -30 -157
rect 30 157 118 170
rect 30 -157 59 157
rect 105 -157 118 157
rect 30 -170 118 -157
rect 184 157 272 170
rect 184 -157 197 157
rect 243 -157 272 157
rect 184 -170 272 -157
rect 332 157 420 170
rect 332 -157 361 157
rect 407 -157 420 157
rect 332 -170 420 -157
rect 486 157 574 170
rect 486 -157 499 157
rect 545 -157 574 157
rect 486 -170 574 -157
rect 634 157 722 170
rect 634 -157 663 157
rect 709 -157 722 157
rect 634 -170 722 -157
rect 788 157 876 170
rect 788 -157 801 157
rect 847 -157 876 157
rect 788 -170 876 -157
rect 936 157 1024 170
rect 936 -157 965 157
rect 1011 -157 1024 157
rect 936 -170 1024 -157
rect 1090 157 1178 170
rect 1090 -157 1103 157
rect 1149 -157 1178 157
rect 1090 -170 1178 -157
rect 1238 157 1326 170
rect 1238 -157 1267 157
rect 1313 -157 1326 157
rect 1238 -170 1326 -157
rect 1392 157 1480 170
rect 1392 -157 1405 157
rect 1451 -157 1480 157
rect 1392 -170 1480 -157
rect 1540 157 1628 170
rect 1540 -157 1569 157
rect 1615 -157 1628 157
rect 1540 -170 1628 -157
rect 1694 157 1782 170
rect 1694 -157 1707 157
rect 1753 -157 1782 157
rect 1694 -170 1782 -157
rect 1842 157 1930 170
rect 1842 -157 1871 157
rect 1917 -157 1930 157
rect 1842 -170 1930 -157
rect 1996 157 2084 170
rect 1996 -157 2009 157
rect 2055 -157 2084 157
rect 1996 -170 2084 -157
rect 2144 157 2232 170
rect 2144 -157 2173 157
rect 2219 -157 2232 157
rect 2144 -170 2232 -157
rect 2298 157 2386 170
rect 2298 -157 2311 157
rect 2357 -157 2386 157
rect 2298 -170 2386 -157
rect 2446 157 2534 170
rect 2446 -157 2475 157
rect 2521 -157 2534 157
rect 2446 -170 2534 -157
<< pdiffc >>
rect -2521 -157 -2475 157
rect -2357 -157 -2311 157
rect -2219 -157 -2173 157
rect -2055 -157 -2009 157
rect -1917 -157 -1871 157
rect -1753 -157 -1707 157
rect -1615 -157 -1569 157
rect -1451 -157 -1405 157
rect -1313 -157 -1267 157
rect -1149 -157 -1103 157
rect -1011 -157 -965 157
rect -847 -157 -801 157
rect -709 -157 -663 157
rect -545 -157 -499 157
rect -407 -157 -361 157
rect -243 -157 -197 157
rect -105 -157 -59 157
rect 59 -157 105 157
rect 197 -157 243 157
rect 361 -157 407 157
rect 499 -157 545 157
rect 663 -157 709 157
rect 801 -157 847 157
rect 965 -157 1011 157
rect 1103 -157 1149 157
rect 1267 -157 1313 157
rect 1405 -157 1451 157
rect 1569 -157 1615 157
rect 1707 -157 1753 157
rect 1871 -157 1917 157
rect 2009 -157 2055 157
rect 2173 -157 2219 157
rect 2311 -157 2357 157
rect 2475 -157 2521 157
<< polysilicon >>
rect -2446 170 -2386 214
rect -2144 170 -2084 214
rect -1842 170 -1782 214
rect -1540 170 -1480 214
rect -1238 170 -1178 214
rect -936 170 -876 214
rect -634 170 -574 214
rect -332 170 -272 214
rect -30 170 30 214
rect 272 170 332 214
rect 574 170 634 214
rect 876 170 936 214
rect 1178 170 1238 214
rect 1480 170 1540 214
rect 1782 170 1842 214
rect 2084 170 2144 214
rect 2386 170 2446 214
rect -2446 -214 -2386 -170
rect -2144 -214 -2084 -170
rect -1842 -214 -1782 -170
rect -1540 -214 -1480 -170
rect -1238 -214 -1178 -170
rect -936 -214 -876 -170
rect -634 -214 -574 -170
rect -332 -214 -272 -170
rect -30 -214 30 -170
rect 272 -214 332 -170
rect 574 -214 634 -170
rect 876 -214 936 -170
rect 1178 -214 1238 -170
rect 1480 -214 1540 -170
rect 1782 -214 1842 -170
rect 2084 -214 2144 -170
rect 2386 -214 2446 -170
<< metal1 >>
rect -2521 157 -2475 168
rect -2521 -168 -2475 -157
rect -2357 157 -2311 168
rect -2357 -168 -2311 -157
rect -2219 157 -2173 168
rect -2219 -168 -2173 -157
rect -2055 157 -2009 168
rect -2055 -168 -2009 -157
rect -1917 157 -1871 168
rect -1917 -168 -1871 -157
rect -1753 157 -1707 168
rect -1753 -168 -1707 -157
rect -1615 157 -1569 168
rect -1615 -168 -1569 -157
rect -1451 157 -1405 168
rect -1451 -168 -1405 -157
rect -1313 157 -1267 168
rect -1313 -168 -1267 -157
rect -1149 157 -1103 168
rect -1149 -168 -1103 -157
rect -1011 157 -965 168
rect -1011 -168 -965 -157
rect -847 157 -801 168
rect -847 -168 -801 -157
rect -709 157 -663 168
rect -709 -168 -663 -157
rect -545 157 -499 168
rect -545 -168 -499 -157
rect -407 157 -361 168
rect -407 -168 -361 -157
rect -243 157 -197 168
rect -243 -168 -197 -157
rect -105 157 -59 168
rect -105 -168 -59 -157
rect 59 157 105 168
rect 59 -168 105 -157
rect 197 157 243 168
rect 197 -168 243 -157
rect 361 157 407 168
rect 361 -168 407 -157
rect 499 157 545 168
rect 499 -168 545 -157
rect 663 157 709 168
rect 663 -168 709 -157
rect 801 157 847 168
rect 801 -168 847 -157
rect 965 157 1011 168
rect 965 -168 1011 -157
rect 1103 157 1149 168
rect 1103 -168 1149 -157
rect 1267 157 1313 168
rect 1267 -168 1313 -157
rect 1405 157 1451 168
rect 1405 -168 1451 -157
rect 1569 157 1615 168
rect 1569 -168 1615 -157
rect 1707 157 1753 168
rect 1707 -168 1753 -157
rect 1871 157 1917 168
rect 1871 -168 1917 -157
rect 2009 157 2055 168
rect 2009 -168 2055 -157
rect 2173 157 2219 168
rect 2173 -168 2219 -157
rect 2311 157 2357 168
rect 2311 -168 2357 -157
rect 2475 157 2521 168
rect 2475 -168 2521 -157
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 1.7 l 0.3 m 1 nf 17 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1757033402
<< nwell >>
rect 330 300 1510 1020
<< pwell >>
rect 330 -250 1510 300
<< nmos >>
rect 580 -30 640 140
rect 770 -30 830 140
rect 1250 -30 1310 140
<< pmos >>
rect 580 460 640 800
rect 770 460 830 800
rect 1250 460 1310 800
<< ndiff >>
rect 459 78 580 140
rect 459 32 492 78
rect 538 32 580 78
rect 459 -30 580 32
rect 640 78 770 140
rect 640 32 682 78
rect 728 32 770 78
rect 640 -30 770 32
rect 830 78 960 140
rect 830 32 872 78
rect 918 32 960 78
rect 1120 78 1250 140
rect 830 -30 960 32
rect 1120 32 1162 78
rect 1208 32 1250 78
rect 1120 -30 1250 32
rect 1310 78 1420 140
rect 1310 32 1352 78
rect 1398 32 1420 78
rect 1310 -30 1420 32
<< pdiff >>
rect 459 563 580 800
rect 459 517 492 563
rect 538 517 580 563
rect 459 460 580 517
rect 640 743 770 800
rect 640 697 682 743
rect 728 697 770 743
rect 640 563 770 697
rect 640 517 682 563
rect 728 517 770 563
rect 640 460 770 517
rect 830 743 960 800
rect 830 697 872 743
rect 918 697 960 743
rect 1120 743 1250 800
rect 830 563 960 697
rect 830 517 872 563
rect 918 517 960 563
rect 830 460 960 517
rect 1120 697 1162 743
rect 1208 697 1250 743
rect 1120 563 1250 697
rect 1120 517 1162 563
rect 1208 517 1250 563
rect 1120 460 1250 517
rect 1310 743 1420 800
rect 1310 697 1352 743
rect 1398 697 1420 743
rect 1310 563 1420 697
rect 1310 517 1352 563
rect 1398 517 1420 563
rect 1310 460 1420 517
<< ndiffc >>
rect 492 32 538 78
rect 682 32 728 78
rect 872 32 918 78
rect 1162 32 1208 78
rect 1352 32 1398 78
<< pdiffc >>
rect 492 517 538 563
rect 682 697 728 743
rect 682 517 728 563
rect 872 697 918 743
rect 872 517 918 563
rect 1162 697 1208 743
rect 1162 517 1208 563
rect 1352 697 1398 743
rect 1352 517 1398 563
<< polysilicon >>
rect 770 850 1100 900
rect 580 800 640 850
rect 770 800 830 850
rect 1020 797 1100 850
rect 1250 800 1310 850
rect 1020 751 1037 797
rect 1083 751 1100 797
rect 1020 700 1100 751
rect 580 360 640 460
rect 770 410 830 460
rect 580 300 830 360
rect 770 290 830 300
rect 1250 290 1310 460
rect 770 263 1310 290
rect 770 217 1212 263
rect 1258 217 1310 263
rect 770 190 1310 217
rect 580 140 640 190
rect 770 140 830 190
rect 1250 140 1310 190
rect 1020 18 1100 70
rect 1020 -28 1037 18
rect 1083 -28 1100 18
rect 580 -130 640 -30
rect 770 -80 830 -30
rect 1020 -130 1100 -28
rect 1250 -80 1310 -30
rect 580 -190 1100 -130
<< polycontact >>
rect 1037 751 1083 797
rect 1212 217 1258 263
rect 1037 -28 1083 18
<< metal1 >>
rect 330 880 1510 1020
rect 330 743 740 800
rect 330 697 682 743
rect 728 697 740 743
rect 330 670 740 697
rect 480 563 550 620
rect 480 517 492 563
rect 538 517 550 563
rect 480 260 550 517
rect 430 170 550 260
rect 480 78 550 170
rect 480 32 492 78
rect 538 32 550 78
rect 480 -30 550 32
rect 670 563 740 670
rect 670 517 682 563
rect 728 517 740 563
rect 670 78 740 517
rect 860 743 930 800
rect 860 697 872 743
rect 918 697 930 743
rect 860 563 930 697
rect 860 517 872 563
rect 918 517 930 563
rect 860 260 930 517
rect 810 170 930 260
rect 670 32 682 78
rect 728 32 740 78
rect 670 -30 740 32
rect 860 78 930 170
rect 860 32 872 78
rect 918 32 930 78
rect 860 -30 930 32
rect 1020 797 1100 830
rect 1020 751 1037 797
rect 1083 751 1100 797
rect 1020 410 1100 751
rect 1150 743 1220 880
rect 1150 697 1162 743
rect 1208 697 1220 743
rect 1150 563 1220 697
rect 1150 517 1162 563
rect 1208 517 1220 563
rect 1150 460 1220 517
rect 1340 743 1450 800
rect 1340 697 1352 743
rect 1398 697 1450 743
rect 1340 563 1450 697
rect 1340 517 1352 563
rect 1398 517 1450 563
rect 1340 460 1450 517
rect 1390 410 1450 460
rect 1020 330 1450 410
rect 1020 18 1100 330
rect 1160 263 1310 280
rect 1160 217 1212 263
rect 1258 217 1310 263
rect 1160 190 1310 217
rect 1390 140 1450 330
rect 1020 -28 1037 18
rect 1083 -28 1100 18
rect 1020 -60 1100 -28
rect 1150 78 1220 140
rect 1150 32 1162 78
rect 1208 32 1220 78
rect 1150 -110 1220 32
rect 1340 78 1450 140
rect 1340 32 1352 78
rect 1398 32 1450 78
rect 1340 -30 1450 32
rect 330 -250 1510 -110
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1755195943
<< pwell >>
rect -2558 -153 2558 153
<< nmos >>
rect -2446 -85 -2386 85
rect -2144 -85 -2084 85
rect -1842 -85 -1782 85
rect -1540 -85 -1480 85
rect -1238 -85 -1178 85
rect -936 -85 -876 85
rect -634 -85 -574 85
rect -332 -85 -272 85
rect -30 -85 30 85
rect 272 -85 332 85
rect 574 -85 634 85
rect 876 -85 936 85
rect 1178 -85 1238 85
rect 1480 -85 1540 85
rect 1782 -85 1842 85
rect 2084 -85 2144 85
rect 2386 -85 2446 85
<< ndiff >>
rect -2534 72 -2446 85
rect -2534 -72 -2521 72
rect -2475 -72 -2446 72
rect -2534 -85 -2446 -72
rect -2386 72 -2298 85
rect -2386 -72 -2357 72
rect -2311 -72 -2298 72
rect -2386 -85 -2298 -72
rect -2232 72 -2144 85
rect -2232 -72 -2219 72
rect -2173 -72 -2144 72
rect -2232 -85 -2144 -72
rect -2084 72 -1996 85
rect -2084 -72 -2055 72
rect -2009 -72 -1996 72
rect -2084 -85 -1996 -72
rect -1930 72 -1842 85
rect -1930 -72 -1917 72
rect -1871 -72 -1842 72
rect -1930 -85 -1842 -72
rect -1782 72 -1694 85
rect -1782 -72 -1753 72
rect -1707 -72 -1694 72
rect -1782 -85 -1694 -72
rect -1628 72 -1540 85
rect -1628 -72 -1615 72
rect -1569 -72 -1540 72
rect -1628 -85 -1540 -72
rect -1480 72 -1392 85
rect -1480 -72 -1451 72
rect -1405 -72 -1392 72
rect -1480 -85 -1392 -72
rect -1326 72 -1238 85
rect -1326 -72 -1313 72
rect -1267 -72 -1238 72
rect -1326 -85 -1238 -72
rect -1178 72 -1090 85
rect -1178 -72 -1149 72
rect -1103 -72 -1090 72
rect -1178 -85 -1090 -72
rect -1024 72 -936 85
rect -1024 -72 -1011 72
rect -965 -72 -936 72
rect -1024 -85 -936 -72
rect -876 72 -788 85
rect -876 -72 -847 72
rect -801 -72 -788 72
rect -876 -85 -788 -72
rect -722 72 -634 85
rect -722 -72 -709 72
rect -663 -72 -634 72
rect -722 -85 -634 -72
rect -574 72 -486 85
rect -574 -72 -545 72
rect -499 -72 -486 72
rect -574 -85 -486 -72
rect -420 72 -332 85
rect -420 -72 -407 72
rect -361 -72 -332 72
rect -420 -85 -332 -72
rect -272 72 -184 85
rect -272 -72 -243 72
rect -197 -72 -184 72
rect -272 -85 -184 -72
rect -118 72 -30 85
rect -118 -72 -105 72
rect -59 -72 -30 72
rect -118 -85 -30 -72
rect 30 72 118 85
rect 30 -72 59 72
rect 105 -72 118 72
rect 30 -85 118 -72
rect 184 72 272 85
rect 184 -72 197 72
rect 243 -72 272 72
rect 184 -85 272 -72
rect 332 72 420 85
rect 332 -72 361 72
rect 407 -72 420 72
rect 332 -85 420 -72
rect 486 72 574 85
rect 486 -72 499 72
rect 545 -72 574 72
rect 486 -85 574 -72
rect 634 72 722 85
rect 634 -72 663 72
rect 709 -72 722 72
rect 634 -85 722 -72
rect 788 72 876 85
rect 788 -72 801 72
rect 847 -72 876 72
rect 788 -85 876 -72
rect 936 72 1024 85
rect 936 -72 965 72
rect 1011 -72 1024 72
rect 936 -85 1024 -72
rect 1090 72 1178 85
rect 1090 -72 1103 72
rect 1149 -72 1178 72
rect 1090 -85 1178 -72
rect 1238 72 1326 85
rect 1238 -72 1267 72
rect 1313 -72 1326 72
rect 1238 -85 1326 -72
rect 1392 72 1480 85
rect 1392 -72 1405 72
rect 1451 -72 1480 72
rect 1392 -85 1480 -72
rect 1540 72 1628 85
rect 1540 -72 1569 72
rect 1615 -72 1628 72
rect 1540 -85 1628 -72
rect 1694 72 1782 85
rect 1694 -72 1707 72
rect 1753 -72 1782 72
rect 1694 -85 1782 -72
rect 1842 72 1930 85
rect 1842 -72 1871 72
rect 1917 -72 1930 72
rect 1842 -85 1930 -72
rect 1996 72 2084 85
rect 1996 -72 2009 72
rect 2055 -72 2084 72
rect 1996 -85 2084 -72
rect 2144 72 2232 85
rect 2144 -72 2173 72
rect 2219 -72 2232 72
rect 2144 -85 2232 -72
rect 2298 72 2386 85
rect 2298 -72 2311 72
rect 2357 -72 2386 72
rect 2298 -85 2386 -72
rect 2446 72 2534 85
rect 2446 -72 2475 72
rect 2521 -72 2534 72
rect 2446 -85 2534 -72
<< ndiffc >>
rect -2521 -72 -2475 72
rect -2357 -72 -2311 72
rect -2219 -72 -2173 72
rect -2055 -72 -2009 72
rect -1917 -72 -1871 72
rect -1753 -72 -1707 72
rect -1615 -72 -1569 72
rect -1451 -72 -1405 72
rect -1313 -72 -1267 72
rect -1149 -72 -1103 72
rect -1011 -72 -965 72
rect -847 -72 -801 72
rect -709 -72 -663 72
rect -545 -72 -499 72
rect -407 -72 -361 72
rect -243 -72 -197 72
rect -105 -72 -59 72
rect 59 -72 105 72
rect 197 -72 243 72
rect 361 -72 407 72
rect 499 -72 545 72
rect 663 -72 709 72
rect 801 -72 847 72
rect 965 -72 1011 72
rect 1103 -72 1149 72
rect 1267 -72 1313 72
rect 1405 -72 1451 72
rect 1569 -72 1615 72
rect 1707 -72 1753 72
rect 1871 -72 1917 72
rect 2009 -72 2055 72
rect 2173 -72 2219 72
rect 2311 -72 2357 72
rect 2475 -72 2521 72
<< polysilicon >>
rect -2446 85 -2386 129
rect -2144 85 -2084 129
rect -1842 85 -1782 129
rect -1540 85 -1480 129
rect -1238 85 -1178 129
rect -936 85 -876 129
rect -634 85 -574 129
rect -332 85 -272 129
rect -30 85 30 129
rect 272 85 332 129
rect 574 85 634 129
rect 876 85 936 129
rect 1178 85 1238 129
rect 1480 85 1540 129
rect 1782 85 1842 129
rect 2084 85 2144 129
rect 2386 85 2446 129
rect -2446 -129 -2386 -85
rect -2144 -129 -2084 -85
rect -1842 -129 -1782 -85
rect -1540 -129 -1480 -85
rect -1238 -129 -1178 -85
rect -936 -129 -876 -85
rect -634 -129 -574 -85
rect -332 -129 -272 -85
rect -30 -129 30 -85
rect 272 -129 332 -85
rect 574 -129 634 -85
rect 876 -129 936 -85
rect 1178 -129 1238 -85
rect 1480 -129 1540 -85
rect 1782 -129 1842 -85
rect 2084 -129 2144 -85
rect 2386 -129 2446 -85
<< metal1 >>
rect -2521 72 -2475 83
rect -2521 -83 -2475 -72
rect -2357 72 -2311 83
rect -2357 -83 -2311 -72
rect -2219 72 -2173 83
rect -2219 -83 -2173 -72
rect -2055 72 -2009 83
rect -2055 -83 -2009 -72
rect -1917 72 -1871 83
rect -1917 -83 -1871 -72
rect -1753 72 -1707 83
rect -1753 -83 -1707 -72
rect -1615 72 -1569 83
rect -1615 -83 -1569 -72
rect -1451 72 -1405 83
rect -1451 -83 -1405 -72
rect -1313 72 -1267 83
rect -1313 -83 -1267 -72
rect -1149 72 -1103 83
rect -1149 -83 -1103 -72
rect -1011 72 -965 83
rect -1011 -83 -965 -72
rect -847 72 -801 83
rect -847 -83 -801 -72
rect -709 72 -663 83
rect -709 -83 -663 -72
rect -545 72 -499 83
rect -545 -83 -499 -72
rect -407 72 -361 83
rect -407 -83 -361 -72
rect -243 72 -197 83
rect -243 -83 -197 -72
rect -105 72 -59 83
rect -105 -83 -59 -72
rect 59 72 105 83
rect 59 -83 105 -72
rect 197 72 243 83
rect 197 -83 243 -72
rect 361 72 407 83
rect 361 -83 407 -72
rect 499 72 545 83
rect 499 -83 545 -72
rect 663 72 709 83
rect 663 -83 709 -72
rect 801 72 847 83
rect 801 -83 847 -72
rect 965 72 1011 83
rect 965 -83 1011 -72
rect 1103 72 1149 83
rect 1103 -83 1149 -72
rect 1267 72 1313 83
rect 1267 -83 1313 -72
rect 1405 72 1451 83
rect 1405 -83 1451 -72
rect 1569 72 1615 83
rect 1569 -83 1615 -72
rect 1707 72 1753 83
rect 1707 -83 1753 -72
rect 1871 72 1917 83
rect 1871 -83 1917 -72
rect 2009 72 2055 83
rect 2009 -83 2055 -72
rect 2173 72 2219 83
rect 2173 -83 2219 -72
rect 2311 72 2357 83
rect 2311 -83 2357 -72
rect 2475 72 2521 83
rect 2475 -83 2521 -72
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.85 l 0.3 m 1 nf 17 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1756212155
<< error_p >>
rect -202 -23 -191 23
rect -34 -23 -23 23
rect 134 -23 145 23
<< nwell >>
rect -290 -159 290 159
<< pmos >>
rect -112 -22 -56 22
rect 56 -22 112 22
<< pdiff >>
rect -204 23 -132 36
rect -204 -23 -191 23
rect -145 22 -132 23
rect -36 23 36 36
rect -36 22 -23 23
rect -145 -22 -112 22
rect -56 -22 -23 22
rect -145 -23 -132 -22
rect -204 -36 -132 -23
rect -36 -23 -23 -22
rect 23 22 36 23
rect 132 23 204 36
rect 132 22 145 23
rect 23 -22 56 22
rect 112 -22 145 22
rect 23 -23 36 -22
rect -36 -36 36 -23
rect 132 -23 145 -22
rect 191 -23 204 23
rect 132 -36 204 -23
<< pdiffc >>
rect -191 -23 -145 23
rect -23 -23 23 23
rect 145 -23 191 23
<< polysilicon >>
rect -112 22 -56 66
rect -112 -66 -56 -22
rect 56 22 112 66
rect 56 -66 112 -22
<< metal1 >>
rect -202 -23 -191 23
rect -145 -23 -134 23
rect -34 -23 -23 23
rect 23 -23 34 23
rect 134 -23 145 23
rect 191 -23 202 23
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.220 l 0.280 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>

** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/sdffrq.sch
.subckt sdffrq VDD D Q SI SE CLK R VSS
*.PININFO D:I SI:I SE:I VDD:B VSS:B Q:O R:I CLK:I
x1 D SI VDD SE VSS net1 mux_2x1
x2 VDD VSS Q net1 CLK R d_flip_flop_r
.ends

* expanding   symbol:  cells/sdffrq/sch/mux_2x1.sym # of pins=6
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/mux_2x1.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/mux_2x1.sch
.subckt mux_2x1 A B VDD S VSS OUT
*.PININFO VDD:B OUT:O A:I B:I S:I VSS:B
x1 VDD S S_INV VSS inv
x2 VDD TG_OUT net1 VSS inv
x3 VDD net1 OUT VSS inv
x4 VDD S A TG_OUT S_INV VSS mux_tg
x5 VDD S_INV B TG_OUT S VSS mux_tg
.ends


* expanding   symbol:  cells/sdffrq/sch/d_flip_flop_r.sym # of pins=6
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/d_flip_flop_r.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/d_flip_flop_r.sch
.subckt d_flip_flop_r VDD VSS Q D CLK R
*.PININFO D:I VDD:I VSS:I Q:O CLK:I R:I
M1 net1 D VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M2 PROBE[0] CLK_INV net2 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M3 PROBE[0] CLK net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M4 net2 D VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M5 CLK_INV CLK VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M8 CLK_INV CLK VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M13 net3 PROBE[1] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M14 PROBE[0] CLK net4 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M15 PROBE[0] CLK_INV net3 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M16 net4 PROBE[1] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M9 net5 PROBE[1] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M10 PROBE[2] CLK net6 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M11 PROBE[2] CLK_INV net5 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M12 net6 PROBE[1] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M19 net7 PROBE[3] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M20 PROBE[2] CLK_INV net8 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M21 PROBE[2] CLK net7 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M22 net8 PROBE[3] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M23 QN PROBE[3] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M24 QN PROBE[3] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M25 Q QN VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M26 Q QN VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M6 net9 PROBE[0] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M27 PROBE[1] R net9 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M28 PROBE[1] PROBE[0] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M17 net10 PROBE[2] VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M29 PROBE[3] R net10 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M30 PROBE[3] PROBE[2] VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M7 PROBE[1] R VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M18 PROBE[3] R VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends


* expanding   symbol:  cells/sdffrq/sch/inv.sym # of pins=4
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/inv.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/inv.sch
.subckt inv VDD IN OUT VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
M2 OUT IN VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M1 OUT IN VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
.ends


* expanding   symbol:  cells/sdffrq/sch/mux_tg.sym # of pins=6
** sym_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/mux_tg.sym
** sch_path: /foss/designs/voidwalkers-scandff-gf180mcu/designs/cells/sdffrq/sch/mux_tg.sch
.subckt mux_tg VDD P_GATE IN OUT N_GATE VSS
*.PININFO VDD:B VSS:B OUT:O IN:I P_GATE:I N_GATE:I
M1 IN N_GATE OUT VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M2 IN P_GATE OUT VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
.ends


magic
tech gf180mcuD
timestamp 1756565017
<< nwell >>
rect -105 65 261 137
<< pwell >>
rect -105 54 261 65
rect -105 52 196 54
rect 209 52 215 54
rect 228 52 234 54
rect 242 52 261 54
rect -105 10 261 52
<< nmos >>
rect -87 32 -81 49
rect -68 32 -62 49
rect -49 32 -43 49
rect -34 32 -28 49
rect 1 32 7 49
rect 12 32 18 49
rect 31 32 37 49
rect 79 32 85 49
rect 118 32 124 49
rect 137 32 143 49
rect 156 32 162 49
rect 171 32 177 49
rect 190 32 196 49
rect 209 32 215 49
rect 228 32 234 49
<< pmos >>
rect -84 81 -78 115
rect -73 81 -67 115
rect -49 81 -43 115
rect -34 81 -28 115
rect -15 81 -9 115
rect 12 81 18 115
rect 31 81 37 115
rect 79 81 85 115
rect 121 81 127 115
rect 137 81 143 115
rect 156 81 162 115
rect 171 81 177 115
rect 190 81 196 115
rect 209 81 215 115
rect 228 81 234 115
<< ndiff >>
rect -98 47 -87 49
rect -98 34 -96 47
rect -91 34 -87 47
rect -98 32 -87 34
rect -81 47 -68 49
rect -81 34 -78 47
rect -71 34 -68 47
rect -81 32 -68 34
rect -62 45 -49 49
rect -62 34 -58 45
rect -53 34 -49 45
rect -62 32 -49 34
rect -43 32 -34 49
rect -28 41 1 49
rect -28 34 -24 41
rect -19 34 1 41
rect -28 32 1 34
rect 7 32 12 49
rect 18 40 31 49
rect 18 34 22 40
rect 27 34 31 40
rect 18 32 31 34
rect 37 47 55 49
rect 37 34 41 47
rect 46 34 55 47
rect 37 32 55 34
rect 68 47 79 49
rect 68 34 70 47
rect 75 34 79 47
rect 68 32 79 34
rect 85 47 100 49
rect 85 34 93 47
rect 98 34 100 47
rect 85 32 100 34
rect 107 47 118 49
rect 107 34 109 47
rect 114 34 118 47
rect 107 32 118 34
rect 124 47 137 49
rect 124 34 127 47
rect 134 34 137 47
rect 124 32 137 34
rect 143 47 156 49
rect 143 34 147 47
rect 152 34 156 47
rect 143 32 156 34
rect 162 32 171 49
rect 177 47 190 49
rect 177 34 181 47
rect 186 34 190 47
rect 177 32 190 34
rect 196 32 209 49
rect 215 47 228 49
rect 215 34 219 47
rect 224 34 228 47
rect 215 32 228 34
rect 234 47 252 49
rect 234 34 238 47
rect 243 34 252 47
rect 234 32 252 34
<< pdiff >>
rect -95 113 -84 115
rect -95 101 -93 113
rect -88 101 -84 113
rect -95 95 -84 101
rect -95 83 -93 95
rect -88 83 -84 95
rect -95 81 -84 83
rect -78 81 -73 115
rect -67 113 -49 115
rect -67 101 -61 113
rect -56 101 -49 113
rect -67 81 -49 101
rect -43 81 -34 115
rect -28 113 -15 115
rect -28 101 -25 113
rect -20 101 -15 113
rect -28 81 -15 101
rect -9 81 12 115
rect 18 113 31 115
rect 18 101 22 113
rect 27 101 31 113
rect 18 81 31 101
rect 37 95 55 115
rect 37 83 46 95
rect 51 83 55 95
rect 37 81 55 83
rect 68 113 79 115
rect 68 101 70 113
rect 75 101 79 113
rect 68 81 79 101
rect 85 95 100 115
rect 85 83 93 95
rect 98 83 100 95
rect 85 81 100 83
rect 110 113 121 115
rect 110 101 112 113
rect 117 101 121 113
rect 110 95 121 101
rect 110 83 112 95
rect 117 83 121 95
rect 110 81 121 83
rect 127 81 137 115
rect 143 113 156 115
rect 143 101 147 113
rect 152 101 156 113
rect 143 95 156 101
rect 143 83 147 95
rect 152 83 156 95
rect 143 81 156 83
rect 162 81 171 115
rect 177 113 190 115
rect 177 101 181 113
rect 186 101 190 113
rect 177 95 190 101
rect 177 83 181 95
rect 186 83 190 95
rect 177 81 190 83
rect 196 81 209 115
rect 215 113 228 115
rect 215 101 219 113
rect 224 101 228 113
rect 215 95 228 101
rect 215 83 219 95
rect 224 83 228 95
rect 215 81 228 83
rect 234 95 252 115
rect 234 83 243 95
rect 248 83 252 95
rect 234 81 252 83
<< ndiffc >>
rect -96 34 -91 47
rect -78 34 -71 47
rect -58 34 -53 45
rect -24 34 -19 41
rect 22 34 27 40
rect 41 34 46 47
rect 70 34 75 47
rect 93 34 98 47
rect 109 34 114 47
rect 127 34 134 47
rect 147 34 152 47
rect 181 34 186 47
rect 219 34 224 47
rect 238 34 243 47
<< pdiffc >>
rect -93 101 -88 113
rect -93 83 -88 95
rect -61 101 -56 113
rect -25 101 -20 113
rect 22 101 27 113
rect 46 83 51 95
rect 70 101 75 113
rect 93 83 98 95
rect 112 101 117 113
rect 112 83 117 95
rect 147 101 152 113
rect 147 83 152 95
rect 181 101 186 113
rect 181 83 186 95
rect 219 101 224 113
rect 219 83 224 95
rect 243 83 248 95
<< polysilicon >>
rect -84 125 85 131
rect -84 115 -78 125
rect -73 115 -67 120
rect -49 115 -43 120
rect -34 115 -28 120
rect -15 115 -9 120
rect 12 115 18 120
rect 31 115 37 120
rect 79 115 85 125
rect 190 125 234 131
rect 121 115 127 120
rect 137 115 143 120
rect 156 115 162 120
rect 171 115 177 120
rect 190 115 196 125
rect 209 115 215 120
rect 228 115 234 125
rect -84 78 -78 81
rect -87 66 -78 78
rect -73 78 -67 81
rect -49 78 -43 81
rect -73 76 -62 78
rect -73 69 -71 76
rect -64 69 -62 76
rect -73 67 -62 69
rect -56 72 -43 78
rect -34 78 -28 81
rect -34 76 -24 78
rect -15 76 -9 81
rect 12 78 18 81
rect 12 76 24 78
rect -87 49 -81 66
rect -73 58 -67 67
rect -56 61 -49 72
rect -34 68 -32 76
rect -26 68 -24 76
rect -34 66 -24 68
rect -17 74 -7 76
rect -17 65 -15 74
rect -9 65 -7 74
rect -17 63 -7 65
rect -2 74 7 76
rect -2 67 0 74
rect 5 67 7 74
rect -56 59 -43 61
rect -73 52 -62 58
rect -56 54 -54 59
rect -49 54 -43 59
rect -15 58 -9 63
rect -56 52 -43 54
rect -68 49 -62 52
rect -49 49 -43 52
rect -34 52 -9 58
rect -2 54 7 67
rect -34 49 -28 52
rect 1 49 7 54
rect 12 70 14 76
rect 22 70 24 76
rect 12 68 24 70
rect 12 49 18 68
rect 31 49 37 81
rect 79 49 85 81
rect 121 78 127 81
rect 111 76 127 78
rect 111 68 113 76
rect 122 68 127 76
rect 111 66 127 68
rect 137 78 143 81
rect 137 76 151 78
rect 137 69 142 76
rect 149 69 151 76
rect 137 67 151 69
rect 118 49 124 66
rect 137 49 143 67
rect 156 65 162 81
rect 171 71 177 81
rect 190 76 196 81
rect 209 78 215 81
rect 209 76 221 78
rect 171 65 196 71
rect 156 63 166 65
rect 156 56 158 63
rect 164 56 166 63
rect 156 54 166 56
rect 190 63 196 65
rect 209 70 211 76
rect 219 70 221 76
rect 209 68 221 70
rect 228 70 234 81
rect 190 61 202 63
rect 190 56 192 61
rect 200 56 202 61
rect 190 54 202 56
rect 156 49 162 54
rect 171 49 177 54
rect 190 49 196 54
rect 209 49 215 68
rect 228 64 258 70
rect 228 49 234 64
rect -87 27 -81 32
rect -68 27 -62 32
rect -49 27 -43 32
rect -34 27 -28 32
rect 1 22 7 32
rect 12 27 18 32
rect 31 22 37 32
rect 79 27 85 32
rect 118 27 124 32
rect 137 27 143 32
rect 156 27 162 32
rect 171 22 177 32
rect 190 27 196 32
rect 209 27 215 32
rect 228 22 234 32
rect 1 16 234 22
<< polycontact >>
rect -71 69 -64 76
rect -32 68 -26 76
rect -15 65 -9 74
rect 0 67 5 74
rect -54 54 -49 59
rect 14 70 22 76
rect 113 68 122 76
rect 142 69 149 76
rect 158 56 164 63
rect 211 70 219 76
rect 192 56 200 61
<< metal1 >>
rect -105 125 261 137
rect -105 113 -87 115
rect -105 102 -93 113
rect -94 101 -93 102
rect -88 101 -87 113
rect -94 95 -87 101
rect -62 113 -55 125
rect -62 101 -61 113
rect -56 101 -55 113
rect -62 99 -55 101
rect -50 113 -18 115
rect -50 101 -25 113
rect -20 101 -18 113
rect -50 99 -18 101
rect 21 113 28 125
rect 21 101 22 113
rect 27 101 28 113
rect 21 99 28 101
rect 33 102 64 115
rect -94 83 -93 95
rect -88 83 -87 95
rect -50 94 -44 99
rect 33 94 40 102
rect -94 61 -87 83
rect -73 88 -44 94
rect -73 76 -62 88
rect -73 69 -71 76
rect -64 72 -62 76
rect -34 82 7 94
rect -34 76 -24 82
rect -64 69 -39 72
rect -73 66 -39 69
rect -34 68 -32 76
rect -26 68 -24 76
rect -34 66 -24 68
rect -15 74 -7 76
rect -94 59 -49 61
rect -94 54 -54 59
rect -78 52 -49 54
rect -97 47 -90 49
rect -97 34 -96 47
rect -91 34 -90 47
rect -97 22 -90 34
rect -78 47 -70 52
rect -71 34 -70 47
rect -78 32 -70 34
rect -59 45 -52 47
rect -59 34 -58 45
rect -53 34 -52 45
rect -59 22 -52 34
rect -44 43 -39 66
rect -9 65 -7 74
rect -15 53 -7 65
rect 0 74 7 82
rect 5 67 7 74
rect 12 88 40 94
rect 45 95 52 97
rect 12 76 24 88
rect 12 70 14 76
rect 22 70 24 76
rect 45 83 46 95
rect 51 83 52 95
rect 57 94 64 102
rect 69 113 76 125
rect 69 101 70 113
rect 75 101 76 113
rect 69 99 76 101
rect 81 113 135 115
rect 81 102 112 113
rect 81 94 87 102
rect 111 101 112 102
rect 117 103 135 113
rect 117 101 118 103
rect 57 87 87 94
rect 92 95 106 97
rect 0 58 7 67
rect 45 53 52 83
rect 92 83 93 95
rect 98 83 106 95
rect 92 81 106 83
rect 111 95 118 101
rect 111 83 112 95
rect 117 83 118 95
rect 111 81 118 83
rect 100 76 106 81
rect 100 68 113 76
rect 122 68 124 76
rect 100 61 106 68
rect -15 47 52 53
rect 92 54 106 61
rect 129 63 135 103
rect 146 113 153 125
rect 146 101 147 113
rect 152 101 153 113
rect 146 95 153 101
rect 146 83 147 95
rect 152 83 153 95
rect 146 81 153 83
rect 158 113 187 115
rect 158 103 181 113
rect 158 76 165 103
rect 140 69 142 76
rect 149 69 165 76
rect 140 68 165 69
rect 180 101 181 103
rect 186 101 187 113
rect 180 95 187 101
rect 180 83 181 95
rect 186 83 187 95
rect 129 56 158 63
rect 164 56 166 63
rect 129 54 166 56
rect -44 41 -18 43
rect -44 34 -24 41
rect -19 34 -18 41
rect -44 32 -18 34
rect 21 40 28 42
rect 21 34 22 40
rect 27 34 28 40
rect 21 22 28 34
rect 40 34 41 47
rect 46 34 52 47
rect 40 32 52 34
rect 69 47 76 49
rect 69 34 70 47
rect 75 34 76 47
rect 69 22 76 34
rect 92 47 99 54
rect 129 49 135 54
rect 92 34 93 47
rect 98 34 99 47
rect 92 32 99 34
rect 108 47 115 49
rect 108 34 109 47
rect 114 34 115 47
rect 108 22 115 34
rect 127 47 135 49
rect 134 34 135 47
rect 127 32 135 34
rect 146 47 153 49
rect 146 34 147 47
rect 152 34 153 47
rect 146 22 153 34
rect 180 47 187 83
rect 218 113 225 125
rect 218 101 219 113
rect 224 101 225 113
rect 218 95 225 101
rect 218 83 219 95
rect 224 83 225 95
rect 218 81 225 83
rect 230 102 252 115
rect 230 76 237 102
rect 209 70 211 76
rect 219 70 237 76
rect 242 95 249 97
rect 242 83 243 95
rect 248 83 249 95
rect 242 63 249 83
rect 192 61 249 63
rect 200 56 249 61
rect 192 54 249 56
rect 242 49 249 54
rect 180 34 181 47
rect 186 34 187 47
rect 180 32 187 34
rect 218 47 225 49
rect 218 34 219 47
rect 224 34 225 47
rect 218 22 225 34
rect 237 47 249 49
rect 237 34 238 47
rect 243 34 249 47
rect 237 32 249 34
rect -105 10 261 22
<< end >>
